typedef enum {RED, GREEN, BLUE, WHITE, ORANGE, CYAN, MAGENTA } LED_COLOR;