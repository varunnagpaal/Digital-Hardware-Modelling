module [module_name]
  /* Parameters Start */
  /* Parameters End */
  /* Port Interface Start */
  /* Port Interface End */
  /* Architecture Start */
    /* Parameter declaration */
    /* Signal declaration */
    /* Component declaration */
    /* Combinational Logic */
    /* Sequential Logic */
  /* Architecture End */
endmodule