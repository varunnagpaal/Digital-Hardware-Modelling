typedef logic unsigned [23:0] color;