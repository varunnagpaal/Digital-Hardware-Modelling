
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_fir_generic_transposed_filter is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_fir_generic_transposed_filter;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_fir_generic_transposed_filter.all;

entity fir_generic_transposed_filter is

   port( clk, rst, valid_x_in : in std_logic;  ready_x_out : out std_logic;  
         valid_h_in : in std_logic;  ready_h_out, valid_out : out std_logic;  
         ready_in : in std_logic;  x_data_in, h_data_in : in SIGNED (15 downto 
         0);  y_data_out : out SIGNED (32 downto 0));

end fir_generic_transposed_filter;

architecture SYN_fir_rtl_arch of fir_generic_transposed_filter is

   component inv
      port( inb : in std_logic;  outb : out std_logic);
   end component;
   
   component xor2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component nand2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component oai22
      port( a, b, c, d : in std_logic;  outb : out std_logic);
   end component;
   
   component aoi22
      port( a, b, c, d : in std_logic;  outb : out std_logic);
   end component;
   
   component nor2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component oai12
      port( b, c, a : in std_logic;  outb : out std_logic);
   end component;
   
   component aoi12
      port( b, c, a : in std_logic;  outb : out std_logic);
   end component;
   
   component dff
      port( d, gclk, rnot : in std_logic;  q : out std_logic);
   end component;
   
   component dff_asyncprehh
      port( d, gclk, asyncprehh : in std_logic;  q : out std_logic);
   end component;
   
   component dff_asyncrsthl
      port( d, gclk, asyncrsthl : in std_logic;  q : out std_logic);
   end component;
   
   signal ready_x_out_port, ready_h_out_port, valid_out_port, 
      coefficient_mem_array_0_15_port, coefficient_mem_array_0_14_port, 
      coefficient_mem_array_0_13_port, coefficient_mem_array_0_12_port, 
      coefficient_mem_array_0_11_port, coefficient_mem_array_0_10_port, 
      coefficient_mem_array_0_9_port, coefficient_mem_array_0_8_port, 
      coefficient_mem_array_0_7_port, coefficient_mem_array_0_6_port, 
      coefficient_mem_array_0_5_port, coefficient_mem_array_0_4_port, 
      coefficient_mem_array_0_3_port, coefficient_mem_array_0_2_port, 
      coefficient_mem_array_0_1_port, coefficient_mem_array_0_0_port, 
      coefficient_mem_array_1_15_port, coefficient_mem_array_1_14_port, 
      coefficient_mem_array_1_13_port, coefficient_mem_array_1_12_port, 
      coefficient_mem_array_1_11_port, coefficient_mem_array_1_10_port, 
      coefficient_mem_array_1_9_port, coefficient_mem_array_1_8_port, 
      coefficient_mem_array_1_7_port, coefficient_mem_array_1_6_port, 
      coefficient_mem_array_1_5_port, coefficient_mem_array_1_4_port, 
      coefficient_mem_array_1_3_port, coefficient_mem_array_1_2_port, 
      coefficient_mem_array_1_1_port, coefficient_mem_array_1_0_port, 
      coefficient_mem_array_2_15_port, coefficient_mem_array_2_14_port, 
      coefficient_mem_array_2_13_port, coefficient_mem_array_2_12_port, 
      coefficient_mem_array_2_11_port, coefficient_mem_array_2_10_port, 
      coefficient_mem_array_2_9_port, coefficient_mem_array_2_8_port, 
      coefficient_mem_array_2_7_port, coefficient_mem_array_2_6_port, 
      coefficient_mem_array_2_5_port, coefficient_mem_array_2_4_port, 
      coefficient_mem_array_2_3_port, coefficient_mem_array_2_2_port, 
      coefficient_mem_array_2_1_port, coefficient_mem_array_2_0_port, 
      coefficient_mem_array_3_15_port, coefficient_mem_array_3_14_port, 
      coefficient_mem_array_3_13_port, coefficient_mem_array_3_12_port, 
      coefficient_mem_array_3_11_port, coefficient_mem_array_3_10_port, 
      coefficient_mem_array_3_9_port, coefficient_mem_array_3_8_port, 
      coefficient_mem_array_3_7_port, coefficient_mem_array_3_6_port, 
      coefficient_mem_array_3_5_port, coefficient_mem_array_3_4_port, 
      coefficient_mem_array_3_3_port, coefficient_mem_array_3_2_port, 
      coefficient_mem_array_3_1_port, coefficient_mem_array_3_0_port, 
      input_sample_mem_15_port, input_sample_mem_14_port, 
      input_sample_mem_13_port, input_sample_mem_12_port, 
      input_sample_mem_11_port, input_sample_mem_10_port, 
      input_sample_mem_9_port, input_sample_mem_8_port, input_sample_mem_7_port
      , input_sample_mem_6_port, input_sample_mem_5_port, 
      input_sample_mem_4_port, input_sample_mem_3_port, input_sample_mem_2_port
      , input_sample_mem_1_port, input_sample_mem_0_port, 
      adder_mem_array_0_32_port, adder_mem_array_0_31_port, 
      adder_mem_array_0_30_port, adder_mem_array_0_29_port, 
      adder_mem_array_0_28_port, adder_mem_array_0_27_port, 
      adder_mem_array_0_26_port, adder_mem_array_0_25_port, 
      adder_mem_array_0_24_port, adder_mem_array_0_23_port, 
      adder_mem_array_0_22_port, adder_mem_array_0_21_port, 
      adder_mem_array_0_20_port, adder_mem_array_0_19_port, 
      adder_mem_array_0_18_port, adder_mem_array_0_17_port, 
      adder_mem_array_0_16_port, adder_mem_array_0_15_port, 
      adder_mem_array_0_14_port, adder_mem_array_0_13_port, 
      adder_mem_array_0_12_port, adder_mem_array_0_11_port, 
      adder_mem_array_0_10_port, adder_mem_array_0_9_port, 
      adder_mem_array_0_8_port, adder_mem_array_0_7_port, 
      adder_mem_array_0_6_port, adder_mem_array_0_5_port, 
      adder_mem_array_0_4_port, adder_mem_array_0_3_port, 
      adder_mem_array_0_2_port, adder_mem_array_0_1_port, 
      adder_mem_array_0_0_port, adder_mem_array_1_32_port, 
      adder_mem_array_1_31_port, adder_mem_array_1_30_port, 
      adder_mem_array_1_29_port, adder_mem_array_1_28_port, 
      adder_mem_array_1_27_port, adder_mem_array_1_26_port, 
      adder_mem_array_1_25_port, adder_mem_array_1_24_port, 
      adder_mem_array_1_23_port, adder_mem_array_1_22_port, 
      adder_mem_array_1_21_port, adder_mem_array_1_20_port, 
      adder_mem_array_1_19_port, adder_mem_array_1_18_port, 
      adder_mem_array_1_17_port, adder_mem_array_1_16_port, 
      adder_mem_array_1_15_port, adder_mem_array_1_14_port, 
      adder_mem_array_1_13_port, adder_mem_array_1_12_port, 
      adder_mem_array_1_11_port, adder_mem_array_1_10_port, 
      adder_mem_array_1_9_port, adder_mem_array_1_8_port, 
      adder_mem_array_1_7_port, adder_mem_array_1_6_port, 
      adder_mem_array_1_5_port, adder_mem_array_1_4_port, 
      adder_mem_array_1_3_port, adder_mem_array_1_2_port, 
      adder_mem_array_1_1_port, adder_mem_array_1_0_port, 
      adder_mem_array_2_32_port, adder_mem_array_2_31_port, 
      adder_mem_array_2_30_port, adder_mem_array_2_29_port, 
      adder_mem_array_2_28_port, adder_mem_array_2_27_port, 
      adder_mem_array_2_26_port, adder_mem_array_2_25_port, 
      adder_mem_array_2_24_port, adder_mem_array_2_23_port, 
      adder_mem_array_2_22_port, adder_mem_array_2_21_port, 
      adder_mem_array_2_20_port, adder_mem_array_2_19_port, 
      adder_mem_array_2_18_port, adder_mem_array_2_17_port, 
      adder_mem_array_2_16_port, adder_mem_array_2_15_port, 
      adder_mem_array_2_14_port, adder_mem_array_2_13_port, 
      adder_mem_array_2_12_port, adder_mem_array_2_11_port, 
      adder_mem_array_2_10_port, adder_mem_array_2_9_port, 
      adder_mem_array_2_8_port, adder_mem_array_2_7_port, 
      adder_mem_array_2_6_port, adder_mem_array_2_5_port, 
      adder_mem_array_2_4_port, adder_mem_array_2_3_port, 
      adder_mem_array_2_2_port, adder_mem_array_2_1_port, 
      adder_mem_array_2_0_port, adder_mem_array_3_32_port, 
      adder_mem_array_3_31_port, adder_mem_array_3_30_port, 
      adder_mem_array_3_29_port, adder_mem_array_3_28_port, 
      adder_mem_array_3_27_port, adder_mem_array_3_26_port, 
      adder_mem_array_3_25_port, adder_mem_array_3_24_port, 
      adder_mem_array_3_23_port, adder_mem_array_3_22_port, 
      adder_mem_array_3_21_port, adder_mem_array_3_20_port, 
      adder_mem_array_3_19_port, adder_mem_array_3_18_port, 
      adder_mem_array_3_17_port, adder_mem_array_3_16_port, 
      adder_mem_array_3_15_port, adder_mem_array_3_14_port, 
      adder_mem_array_3_13_port, adder_mem_array_3_12_port, 
      adder_mem_array_3_11_port, adder_mem_array_3_10_port, 
      adder_mem_array_3_9_port, adder_mem_array_3_8_port, 
      adder_mem_array_3_7_port, adder_mem_array_3_6_port, 
      adder_mem_array_3_5_port, adder_mem_array_3_4_port, 
      adder_mem_array_3_3_port, adder_mem_array_3_2_port, 
      adder_mem_array_3_1_port, adder_mem_array_3_0_port, 
      multiplier_sigs_0_31_port, multiplier_sigs_0_30_port, 
      multiplier_sigs_0_29_port, multiplier_sigs_0_28_port, 
      multiplier_sigs_0_27_port, multiplier_sigs_0_26_port, 
      multiplier_sigs_0_25_port, multiplier_sigs_0_24_port, 
      multiplier_sigs_0_23_port, multiplier_sigs_0_22_port, 
      multiplier_sigs_0_21_port, multiplier_sigs_0_20_port, 
      multiplier_sigs_0_19_port, multiplier_sigs_0_18_port, 
      multiplier_sigs_0_17_port, multiplier_sigs_0_16_port, 
      multiplier_sigs_0_15_port, multiplier_sigs_0_14_port, 
      multiplier_sigs_0_13_port, multiplier_sigs_0_12_port, 
      multiplier_sigs_0_11_port, multiplier_sigs_0_10_port, 
      multiplier_sigs_0_9_port, multiplier_sigs_0_8_port, 
      multiplier_sigs_0_7_port, multiplier_sigs_0_6_port, 
      multiplier_sigs_0_5_port, multiplier_sigs_0_4_port, 
      multiplier_sigs_0_3_port, multiplier_sigs_0_2_port, 
      multiplier_sigs_0_0_port, multiplier_sigs_1_31_port, 
      multiplier_sigs_1_30_port, multiplier_sigs_1_29_port, 
      multiplier_sigs_1_28_port, multiplier_sigs_1_27_port, 
      multiplier_sigs_1_26_port, multiplier_sigs_1_25_port, 
      multiplier_sigs_1_24_port, multiplier_sigs_1_23_port, 
      multiplier_sigs_1_22_port, multiplier_sigs_1_21_port, 
      multiplier_sigs_1_20_port, multiplier_sigs_1_19_port, 
      multiplier_sigs_1_18_port, multiplier_sigs_1_17_port, 
      multiplier_sigs_1_16_port, multiplier_sigs_1_15_port, 
      multiplier_sigs_1_14_port, multiplier_sigs_1_13_port, 
      multiplier_sigs_1_12_port, multiplier_sigs_1_11_port, 
      multiplier_sigs_1_10_port, multiplier_sigs_1_9_port, 
      multiplier_sigs_1_8_port, multiplier_sigs_1_7_port, 
      multiplier_sigs_1_6_port, multiplier_sigs_1_5_port, 
      multiplier_sigs_1_4_port, multiplier_sigs_1_3_port, 
      multiplier_sigs_1_2_port, multiplier_sigs_1_0_port, 
      multiplier_sigs_2_31_port, multiplier_sigs_2_30_port, 
      multiplier_sigs_2_29_port, multiplier_sigs_2_28_port, 
      multiplier_sigs_2_27_port, multiplier_sigs_2_26_port, 
      multiplier_sigs_2_25_port, multiplier_sigs_2_24_port, 
      multiplier_sigs_2_23_port, multiplier_sigs_2_22_port, 
      multiplier_sigs_2_21_port, multiplier_sigs_2_20_port, 
      multiplier_sigs_2_19_port, multiplier_sigs_2_18_port, 
      multiplier_sigs_2_17_port, multiplier_sigs_2_16_port, 
      multiplier_sigs_2_15_port, multiplier_sigs_2_14_port, 
      multiplier_sigs_2_13_port, multiplier_sigs_2_12_port, 
      multiplier_sigs_2_11_port, multiplier_sigs_2_10_port, 
      multiplier_sigs_2_9_port, multiplier_sigs_2_8_port, 
      multiplier_sigs_2_7_port, multiplier_sigs_2_6_port, 
      multiplier_sigs_2_5_port, multiplier_sigs_2_4_port, 
      multiplier_sigs_2_3_port, multiplier_sigs_2_2_port, 
      multiplier_sigs_2_0_port, multiplier_sigs_3_31_port, 
      multiplier_sigs_3_30_port, multiplier_sigs_3_29_port, 
      multiplier_sigs_3_28_port, multiplier_sigs_3_27_port, 
      multiplier_sigs_3_26_port, multiplier_sigs_3_25_port, 
      multiplier_sigs_3_24_port, multiplier_sigs_3_23_port, 
      multiplier_sigs_3_22_port, multiplier_sigs_3_21_port, 
      multiplier_sigs_3_20_port, multiplier_sigs_3_19_port, 
      multiplier_sigs_3_18_port, multiplier_sigs_3_17_port, 
      multiplier_sigs_3_16_port, multiplier_sigs_3_15_port, 
      multiplier_sigs_3_14_port, multiplier_sigs_3_13_port, 
      multiplier_sigs_3_12_port, multiplier_sigs_3_11_port, 
      multiplier_sigs_3_10_port, multiplier_sigs_3_9_port, 
      multiplier_sigs_3_8_port, multiplier_sigs_3_7_port, 
      multiplier_sigs_3_6_port, multiplier_sigs_3_5_port, 
      multiplier_sigs_3_4_port, multiplier_sigs_3_3_port, 
      multiplier_sigs_3_2_port, multiplier_sigs_3_1_port, 
      multiplier_sigs_3_0_port, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, 
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, 
      N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59
      , N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, 
      N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88
      , N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102
      , N103, N104, coeff_cnt_1_port, coeff_cnt_0_port, n16_port, n17_port, 
      n18_port, n19_port, n20_port, n21_port, n22_port, n23_port, n24_port, 
      n25_port, n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, 
      n32_port, n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, 
      n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, 
      n46_port, n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, 
      n53_port, n54_port, n55_port, n56_port, n57_port, n58_port, n59_port, 
      n60_port, n61_port, n62_port, n63_port, n64_port, n65_port, n66_port, 
      n67_port, n68_port, n69_port, n70_port, n71_port, n72_port, n73_port, 
      n74_port, n75_port, n76_port, n77_port, n78_port, n79_port, n80_port, 
      n81_port, n82_port, n83_port, n84_port, n85_port, n86_port, n87_port, 
      n88_port, n89_port, n90_port, n91_port, n92_port, n93_port, n94_port, 
      n95_port, n96_port, n97_port, n98_port, n99_port, n100_port, n101_port, 
      n102_port, n103_port, n104_port, n105, n106, n107, n108, n109, n110, n111
      , n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, 
      mult_125_G3_FS_1_C_1_3_3_port, mult_125_G3_FS_1_C_1_4_0_port, 
      mult_125_G3_FS_1_C_1_4_1_port, mult_125_G3_FS_1_C_1_4_2_port, 
      mult_125_G3_FS_1_C_1_4_3_port, mult_125_G3_FS_1_C_1_5_0_port, 
      mult_125_G3_FS_1_C_1_5_1_port, mult_125_G3_FS_1_C_1_5_2_port, 
      mult_125_G3_FS_1_C_1_5_3_port, mult_125_G3_FS_1_C_1_6_0_port, 
      mult_125_G3_FS_1_C_1_6_1_port, mult_125_G3_FS_1_C_1_6_2_port, 
      mult_125_G3_FS_1_C_1_6_3_port, mult_125_G3_FS_1_C_1_7_0_port, 
      mult_125_G3_FS_1_C_1_7_1_port, mult_125_G3_FS_1_P_0_0_1_port, 
      mult_125_G3_FS_1_P_0_0_2_port, mult_125_G3_FS_1_P_0_0_3_port, 
      mult_125_G3_FS_1_P_0_1_1_port, mult_125_G3_FS_1_P_0_1_2_port, 
      mult_125_G3_FS_1_P_0_1_3_port, mult_125_G3_FS_1_P_0_2_1_port, 
      mult_125_G3_FS_1_P_0_2_2_port, mult_125_G3_FS_1_P_0_2_3_port, 
      mult_125_G3_FS_1_P_0_3_1_port, mult_125_G3_FS_1_P_0_3_2_port, 
      mult_125_G3_FS_1_P_0_3_3_port, mult_125_G3_FS_1_P_0_4_1_port, 
      mult_125_G3_FS_1_P_0_4_2_port, mult_125_G3_FS_1_P_0_4_3_port, 
      mult_125_G3_FS_1_P_0_5_1_port, mult_125_G3_FS_1_P_0_5_2_port, 
      mult_125_G3_FS_1_P_0_5_3_port, mult_125_G3_FS_1_P_0_6_1_port, 
      mult_125_G3_FS_1_P_0_6_2_port, mult_125_G3_FS_1_P_0_6_3_port, 
      mult_125_G3_FS_1_P_0_7_1_port, mult_125_G3_FS_1_TEMP_P_0_0_0_port, 
      mult_125_G3_FS_1_TEMP_P_0_1_0_port, mult_125_G3_FS_1_TEMP_P_0_2_0_port, 
      mult_125_G3_FS_1_TEMP_P_0_3_0_port, mult_125_G3_FS_1_TEMP_P_0_4_0_port, 
      mult_125_G3_FS_1_TEMP_P_0_4_1_port, mult_125_G3_FS_1_TEMP_P_0_4_2_port, 
      mult_125_G3_FS_1_TEMP_P_0_5_0_port, mult_125_G3_FS_1_TEMP_P_0_5_1_port, 
      mult_125_G3_FS_1_TEMP_P_0_5_2_port, mult_125_G3_FS_1_TEMP_P_0_6_0_port, 
      mult_125_G3_FS_1_TEMP_P_0_6_1_port, mult_125_G3_FS_1_TEMP_P_0_6_2_port, 
      mult_125_G3_FS_1_TEMP_P_0_7_0_port, mult_125_G3_FS_1_G_1_0_3_port, 
      mult_125_G3_FS_1_G_1_1_0_port, mult_125_G3_FS_1_G_1_1_1_port, 
      mult_125_G3_FS_1_G_1_1_2_port, mult_125_G3_FS_1_G_2_0_0_port, 
      mult_125_G3_FS_1_TEMP_G_0_3_2_port, mult_125_G3_FS_1_TEMP_G_0_4_1_port, 
      mult_125_G3_FS_1_TEMP_G_0_4_2_port, mult_125_G3_FS_1_TEMP_G_0_5_1_port, 
      mult_125_G3_FS_1_TEMP_G_0_5_2_port, mult_125_G3_FS_1_TEMP_G_0_6_1_port, 
      mult_125_G3_FS_1_TEMP_G_0_6_2_port, mult_125_G3_FS_1_G_n_int_0_3_2_port, 
      mult_125_G3_FS_1_G_n_int_0_3_3_port, mult_125_G3_FS_1_G_n_int_0_4_0_port,
      mult_125_G3_FS_1_G_n_int_0_4_1_port, mult_125_G3_FS_1_G_n_int_0_4_2_port,
      mult_125_G3_FS_1_G_n_int_0_4_3_port, mult_125_G3_FS_1_G_n_int_0_5_0_port,
      mult_125_G3_FS_1_G_n_int_0_5_1_port, mult_125_G3_FS_1_G_n_int_0_5_2_port,
      mult_125_G3_FS_1_G_n_int_0_5_3_port, mult_125_G3_FS_1_G_n_int_0_6_0_port,
      mult_125_G3_FS_1_G_n_int_0_6_1_port, mult_125_G3_FS_1_G_n_int_0_6_2_port,
      mult_125_G3_FS_1_G_n_int_0_6_3_port, mult_125_G3_FS_1_G_n_int_0_7_0_port,
      mult_125_G3_FS_1_G_n_int_0_7_1_port, mult_125_G3_FS_1_PG_int_0_3_3_port, 
      mult_125_G3_FS_1_PG_int_0_4_0_port, mult_125_G3_FS_1_PG_int_0_4_1_port, 
      mult_125_G3_FS_1_PG_int_0_4_2_port, mult_125_G3_FS_1_PG_int_0_4_3_port, 
      mult_125_G3_FS_1_PG_int_0_5_0_port, mult_125_G3_FS_1_PG_int_0_5_1_port, 
      mult_125_G3_FS_1_PG_int_0_5_2_port, mult_125_G3_FS_1_PG_int_0_5_3_port, 
      mult_125_G3_FS_1_PG_int_0_6_0_port, mult_125_G3_FS_1_PG_int_0_6_1_port, 
      mult_125_G3_FS_1_PG_int_0_6_2_port, mult_125_G3_FS_1_PG_int_0_6_3_port, 
      mult_125_G3_FS_1_PG_int_0_7_0_port, mult_125_G3_FS_1_PG_int_0_7_1_port, 
      mult_125_G3_A2_14_port, mult_125_G3_A2_15_port, mult_125_G3_A2_16_port, 
      mult_125_G3_A2_17_port, mult_125_G3_A2_18_port, mult_125_G3_A2_19_port, 
      mult_125_G3_A2_20_port, mult_125_G3_A2_21_port, mult_125_G3_A2_22_port, 
      mult_125_G3_A2_23_port, mult_125_G3_A2_24_port, mult_125_G3_A2_25_port, 
      mult_125_G3_A2_26_port, mult_125_G3_A2_27_port, mult_125_G3_A2_28_port, 
      mult_125_G3_A2_29_port, mult_125_G3_A1_0_port, mult_125_G3_A1_1_port, 
      mult_125_G3_A1_2_port, mult_125_G3_A1_3_port, mult_125_G3_A1_4_port, 
      mult_125_G3_A1_5_port, mult_125_G3_A1_6_port, mult_125_G3_A1_7_port, 
      mult_125_G3_A1_8_port, mult_125_G3_A1_9_port, mult_125_G3_A1_10_port, 
      mult_125_G3_A1_11_port, mult_125_G3_A1_12_port, mult_125_G3_A1_13_port, 
      mult_125_G3_A1_14_port, mult_125_G3_A1_15_port, mult_125_G3_A1_16_port, 
      mult_125_G3_A1_17_port, mult_125_G3_A1_18_port, mult_125_G3_A1_19_port, 
      mult_125_G3_A1_20_port, mult_125_G3_A1_21_port, mult_125_G3_A1_22_port, 
      mult_125_G3_A1_23_port, mult_125_G3_A1_24_port, mult_125_G3_A1_25_port, 
      mult_125_G3_A1_26_port, mult_125_G3_A1_27_port, mult_125_G3_A1_28_port, 
      mult_125_G3_A1_29_port, mult_125_G3_ZB, mult_125_G3_ZA, mult_125_G3_QB, 
      mult_125_G3_QA, mult_125_G3_A_notx_0_port, mult_125_G3_A_notx_1_port, 
      mult_125_G3_A_notx_2_port, mult_125_G3_A_notx_3_port, 
      mult_125_G3_A_notx_4_port, mult_125_G3_A_notx_5_port, 
      mult_125_G3_A_notx_6_port, mult_125_G3_A_notx_7_port, 
      mult_125_G3_A_notx_8_port, mult_125_G3_A_notx_9_port, 
      mult_125_G3_A_notx_10_port, mult_125_G3_A_notx_11_port, 
      mult_125_G3_A_notx_12_port, mult_125_G3_A_notx_13_port, 
      mult_125_G3_A_notx_14_port, mult_125_G3_B_notx_0_port, 
      mult_125_G3_B_notx_1_port, mult_125_G3_B_notx_2_port, 
      mult_125_G3_B_notx_3_port, mult_125_G3_B_notx_4_port, 
      mult_125_G3_B_notx_5_port, mult_125_G3_B_notx_6_port, 
      mult_125_G3_B_notx_7_port, mult_125_G3_B_notx_8_port, 
      mult_125_G3_B_notx_9_port, mult_125_G3_B_notx_10_port, 
      mult_125_G3_B_notx_11_port, mult_125_G3_B_notx_12_port, 
      mult_125_G3_B_notx_13_port, mult_125_G3_B_notx_14_port, 
      mult_125_G3_ab_0_1_port, mult_125_G3_ab_0_2_port, mult_125_G3_ab_0_3_port
      , mult_125_G3_ab_0_4_port, mult_125_G3_ab_0_5_port, 
      mult_125_G3_ab_0_6_port, mult_125_G3_ab_0_7_port, mult_125_G3_ab_0_8_port
      , mult_125_G3_ab_0_9_port, mult_125_G3_ab_0_10_port, 
      mult_125_G3_ab_0_11_port, mult_125_G3_ab_0_12_port, 
      mult_125_G3_ab_0_13_port, mult_125_G3_ab_0_14_port, 
      mult_125_G3_ab_0_15_port, mult_125_G3_ab_1_0_port, 
      mult_125_G3_ab_1_1_port, mult_125_G3_ab_1_2_port, mult_125_G3_ab_1_3_port
      , mult_125_G3_ab_1_4_port, mult_125_G3_ab_1_5_port, 
      mult_125_G3_ab_1_6_port, mult_125_G3_ab_1_7_port, mult_125_G3_ab_1_8_port
      , mult_125_G3_ab_1_9_port, mult_125_G3_ab_1_10_port, 
      mult_125_G3_ab_1_11_port, mult_125_G3_ab_1_12_port, 
      mult_125_G3_ab_1_13_port, mult_125_G3_ab_1_14_port, 
      mult_125_G3_ab_1_15_port, mult_125_G3_ab_2_0_port, 
      mult_125_G3_ab_2_1_port, mult_125_G3_ab_2_2_port, mult_125_G3_ab_2_3_port
      , mult_125_G3_ab_2_4_port, mult_125_G3_ab_2_5_port, 
      mult_125_G3_ab_2_6_port, mult_125_G3_ab_2_7_port, mult_125_G3_ab_2_8_port
      , mult_125_G3_ab_2_9_port, mult_125_G3_ab_2_10_port, 
      mult_125_G3_ab_2_11_port, mult_125_G3_ab_2_12_port, 
      mult_125_G3_ab_2_13_port, mult_125_G3_ab_2_14_port, 
      mult_125_G3_ab_2_15_port, mult_125_G3_ab_3_0_port, 
      mult_125_G3_ab_3_1_port, mult_125_G3_ab_3_2_port, mult_125_G3_ab_3_3_port
      , mult_125_G3_ab_3_4_port, mult_125_G3_ab_3_5_port, 
      mult_125_G3_ab_3_6_port, mult_125_G3_ab_3_7_port, mult_125_G3_ab_3_8_port
      , mult_125_G3_ab_3_9_port, mult_125_G3_ab_3_10_port, 
      mult_125_G3_ab_3_11_port, mult_125_G3_ab_3_12_port, 
      mult_125_G3_ab_3_13_port, mult_125_G3_ab_3_14_port, 
      mult_125_G3_ab_3_15_port, mult_125_G3_ab_4_0_port, 
      mult_125_G3_ab_4_1_port, mult_125_G3_ab_4_2_port, mult_125_G3_ab_4_3_port
      , mult_125_G3_ab_4_4_port, mult_125_G3_ab_4_5_port, 
      mult_125_G3_ab_4_6_port, mult_125_G3_ab_4_7_port, mult_125_G3_ab_4_8_port
      , mult_125_G3_ab_4_9_port, mult_125_G3_ab_4_10_port, 
      mult_125_G3_ab_4_11_port, mult_125_G3_ab_4_12_port, 
      mult_125_G3_ab_4_13_port, mult_125_G3_ab_4_14_port, 
      mult_125_G3_ab_4_15_port, mult_125_G3_ab_5_0_port, 
      mult_125_G3_ab_5_1_port, mult_125_G3_ab_5_2_port, mult_125_G3_ab_5_3_port
      , mult_125_G3_ab_5_4_port, mult_125_G3_ab_5_5_port, 
      mult_125_G3_ab_5_6_port, mult_125_G3_ab_5_7_port, mult_125_G3_ab_5_8_port
      , mult_125_G3_ab_5_9_port, mult_125_G3_ab_5_10_port, 
      mult_125_G3_ab_5_11_port, mult_125_G3_ab_5_12_port, 
      mult_125_G3_ab_5_13_port, mult_125_G3_ab_5_14_port, 
      mult_125_G3_ab_5_15_port, mult_125_G3_ab_6_0_port, 
      mult_125_G3_ab_6_1_port, mult_125_G3_ab_6_2_port, mult_125_G3_ab_6_3_port
      , mult_125_G3_ab_6_4_port, mult_125_G3_ab_6_5_port, 
      mult_125_G3_ab_6_6_port, mult_125_G3_ab_6_7_port, mult_125_G3_ab_6_8_port
      , mult_125_G3_ab_6_9_port, mult_125_G3_ab_6_10_port, 
      mult_125_G3_ab_6_11_port, mult_125_G3_ab_6_12_port, 
      mult_125_G3_ab_6_13_port, mult_125_G3_ab_6_14_port, 
      mult_125_G3_ab_6_15_port, mult_125_G3_ab_7_0_port, 
      mult_125_G3_ab_7_1_port, mult_125_G3_ab_7_2_port, mult_125_G3_ab_7_3_port
      , mult_125_G3_ab_7_4_port, mult_125_G3_ab_7_5_port, 
      mult_125_G3_ab_7_6_port, mult_125_G3_ab_7_7_port, mult_125_G3_ab_7_8_port
      , mult_125_G3_ab_7_9_port, mult_125_G3_ab_7_10_port, 
      mult_125_G3_ab_7_11_port, mult_125_G3_ab_7_12_port, 
      mult_125_G3_ab_7_13_port, mult_125_G3_ab_7_14_port, 
      mult_125_G3_ab_7_15_port, mult_125_G3_ab_8_0_port, 
      mult_125_G3_ab_8_1_port, mult_125_G3_ab_8_2_port, mult_125_G3_ab_8_3_port
      , mult_125_G3_ab_8_4_port, mult_125_G3_ab_8_5_port, 
      mult_125_G3_ab_8_6_port, mult_125_G3_ab_8_7_port, mult_125_G3_ab_8_8_port
      , mult_125_G3_ab_8_9_port, mult_125_G3_ab_8_10_port, 
      mult_125_G3_ab_8_11_port, mult_125_G3_ab_8_12_port, 
      mult_125_G3_ab_8_13_port, mult_125_G3_ab_8_14_port, 
      mult_125_G3_ab_8_15_port, mult_125_G3_ab_9_0_port, 
      mult_125_G3_ab_9_1_port, mult_125_G3_ab_9_2_port, mult_125_G3_ab_9_3_port
      , mult_125_G3_ab_9_4_port, mult_125_G3_ab_9_5_port, 
      mult_125_G3_ab_9_6_port, mult_125_G3_ab_9_7_port, mult_125_G3_ab_9_8_port
      , mult_125_G3_ab_9_9_port, mult_125_G3_ab_9_10_port, 
      mult_125_G3_ab_9_11_port, mult_125_G3_ab_9_12_port, 
      mult_125_G3_ab_9_13_port, mult_125_G3_ab_9_14_port, 
      mult_125_G3_ab_9_15_port, mult_125_G3_ab_10_0_port, 
      mult_125_G3_ab_10_1_port, mult_125_G3_ab_10_2_port, 
      mult_125_G3_ab_10_3_port, mult_125_G3_ab_10_4_port, 
      mult_125_G3_ab_10_5_port, mult_125_G3_ab_10_6_port, 
      mult_125_G3_ab_10_7_port, mult_125_G3_ab_10_8_port, 
      mult_125_G3_ab_10_9_port, mult_125_G3_ab_10_10_port, 
      mult_125_G3_ab_10_11_port, mult_125_G3_ab_10_12_port, 
      mult_125_G3_ab_10_13_port, mult_125_G3_ab_10_14_port, 
      mult_125_G3_ab_10_15_port, mult_125_G3_ab_11_0_port, 
      mult_125_G3_ab_11_1_port, mult_125_G3_ab_11_2_port, 
      mult_125_G3_ab_11_3_port, mult_125_G3_ab_11_4_port, 
      mult_125_G3_ab_11_5_port, mult_125_G3_ab_11_6_port, 
      mult_125_G3_ab_11_7_port, mult_125_G3_ab_11_8_port, 
      mult_125_G3_ab_11_9_port, mult_125_G3_ab_11_10_port, 
      mult_125_G3_ab_11_11_port, mult_125_G3_ab_11_12_port, 
      mult_125_G3_ab_11_13_port, mult_125_G3_ab_11_14_port, 
      mult_125_G3_ab_11_15_port, mult_125_G3_ab_12_0_port, 
      mult_125_G3_ab_12_1_port, mult_125_G3_ab_12_2_port, 
      mult_125_G3_ab_12_3_port, mult_125_G3_ab_12_4_port, 
      mult_125_G3_ab_12_5_port, mult_125_G3_ab_12_6_port, 
      mult_125_G3_ab_12_7_port, mult_125_G3_ab_12_8_port, 
      mult_125_G3_ab_12_9_port, mult_125_G3_ab_12_10_port, 
      mult_125_G3_ab_12_11_port, mult_125_G3_ab_12_12_port, 
      mult_125_G3_ab_12_13_port, mult_125_G3_ab_12_14_port, 
      mult_125_G3_ab_12_15_port, mult_125_G3_ab_13_0_port, 
      mult_125_G3_ab_13_1_port, mult_125_G3_ab_13_2_port, 
      mult_125_G3_ab_13_3_port, mult_125_G3_ab_13_4_port, 
      mult_125_G3_ab_13_5_port, mult_125_G3_ab_13_6_port, 
      mult_125_G3_ab_13_7_port, mult_125_G3_ab_13_8_port, 
      mult_125_G3_ab_13_9_port, mult_125_G3_ab_13_10_port, 
      mult_125_G3_ab_13_11_port, mult_125_G3_ab_13_12_port, 
      mult_125_G3_ab_13_13_port, mult_125_G3_ab_13_14_port, 
      mult_125_G3_ab_13_15_port, mult_125_G3_ab_14_0_port, 
      mult_125_G3_ab_14_1_port, mult_125_G3_ab_14_2_port, 
      mult_125_G3_ab_14_3_port, mult_125_G3_ab_14_4_port, 
      mult_125_G3_ab_14_5_port, mult_125_G3_ab_14_6_port, 
      mult_125_G3_ab_14_7_port, mult_125_G3_ab_14_8_port, 
      mult_125_G3_ab_14_9_port, mult_125_G3_ab_14_10_port, 
      mult_125_G3_ab_14_11_port, mult_125_G3_ab_14_12_port, 
      mult_125_G3_ab_14_13_port, mult_125_G3_ab_14_14_port, 
      mult_125_G3_ab_14_15_port, mult_125_G3_ab_15_0_port, 
      mult_125_G3_ab_15_1_port, mult_125_G3_ab_15_2_port, 
      mult_125_G3_ab_15_3_port, mult_125_G3_ab_15_4_port, 
      mult_125_G3_ab_15_5_port, mult_125_G3_ab_15_6_port, 
      mult_125_G3_ab_15_7_port, mult_125_G3_ab_15_8_port, 
      mult_125_G3_ab_15_9_port, mult_125_G3_ab_15_10_port, 
      mult_125_G3_ab_15_11_port, mult_125_G3_ab_15_12_port, 
      mult_125_G3_ab_15_13_port, mult_125_G3_ab_15_14_port, 
      mult_125_G3_ab_15_15_port, mult_125_G3_B_not_0_port, 
      mult_125_G3_B_not_1_port, mult_125_G3_B_not_2_port, 
      mult_125_G3_B_not_3_port, mult_125_G3_B_not_4_port, 
      mult_125_G3_B_not_5_port, mult_125_G3_B_not_6_port, 
      mult_125_G3_B_not_7_port, mult_125_G3_B_not_8_port, 
      mult_125_G3_B_not_9_port, mult_125_G3_B_not_10_port, 
      mult_125_G3_B_not_11_port, mult_125_G3_B_not_12_port, 
      mult_125_G3_B_not_13_port, mult_125_G3_B_not_14_port, 
      mult_125_G3_B_not_15_port, mult_125_G3_A_not_0_port, 
      mult_125_G3_A_not_1_port, mult_125_G3_A_not_2_port, 
      mult_125_G3_A_not_3_port, mult_125_G3_A_not_4_port, 
      mult_125_G3_A_not_5_port, mult_125_G3_A_not_6_port, 
      mult_125_G3_A_not_7_port, mult_125_G3_A_not_8_port, 
      mult_125_G3_A_not_9_port, mult_125_G3_A_not_10_port, 
      mult_125_G3_A_not_11_port, mult_125_G3_A_not_12_port, 
      mult_125_G3_A_not_13_port, mult_125_G3_A_not_14_port, 
      mult_125_G3_A_not_15_port, mult_125_G2_FS_1_C_1_3_3_port, 
      mult_125_G2_FS_1_C_1_4_0_port, mult_125_G2_FS_1_C_1_4_1_port, 
      mult_125_G2_FS_1_C_1_4_2_port, mult_125_G2_FS_1_C_1_4_3_port, 
      mult_125_G2_FS_1_C_1_5_0_port, mult_125_G2_FS_1_C_1_5_1_port, 
      mult_125_G2_FS_1_C_1_5_2_port, mult_125_G2_FS_1_C_1_5_3_port, 
      mult_125_G2_FS_1_C_1_6_0_port, mult_125_G2_FS_1_C_1_6_1_port, 
      mult_125_G2_FS_1_C_1_6_2_port, mult_125_G2_FS_1_C_1_6_3_port, 
      mult_125_G2_FS_1_C_1_7_0_port, mult_125_G2_FS_1_C_1_7_1_port, 
      mult_125_G2_FS_1_P_0_0_1_port, mult_125_G2_FS_1_P_0_0_2_port, 
      mult_125_G2_FS_1_P_0_0_3_port, mult_125_G2_FS_1_P_0_1_1_port, 
      mult_125_G2_FS_1_P_0_1_2_port, mult_125_G2_FS_1_P_0_1_3_port, 
      mult_125_G2_FS_1_P_0_2_1_port, mult_125_G2_FS_1_P_0_2_2_port, 
      mult_125_G2_FS_1_P_0_2_3_port, mult_125_G2_FS_1_P_0_3_1_port, 
      mult_125_G2_FS_1_P_0_3_2_port, mult_125_G2_FS_1_P_0_3_3_port, 
      mult_125_G2_FS_1_P_0_4_1_port, mult_125_G2_FS_1_P_0_4_2_port, 
      mult_125_G2_FS_1_P_0_4_3_port, mult_125_G2_FS_1_P_0_5_1_port, 
      mult_125_G2_FS_1_P_0_5_2_port, mult_125_G2_FS_1_P_0_5_3_port, 
      mult_125_G2_FS_1_P_0_6_1_port, mult_125_G2_FS_1_P_0_6_2_port, 
      mult_125_G2_FS_1_P_0_6_3_port, mult_125_G2_FS_1_P_0_7_1_port, 
      mult_125_G2_FS_1_TEMP_P_0_0_0_port, mult_125_G2_FS_1_TEMP_P_0_1_0_port, 
      mult_125_G2_FS_1_TEMP_P_0_2_0_port, mult_125_G2_FS_1_TEMP_P_0_3_0_port, 
      mult_125_G2_FS_1_TEMP_P_0_4_0_port, mult_125_G2_FS_1_TEMP_P_0_4_1_port, 
      mult_125_G2_FS_1_TEMP_P_0_4_2_port, mult_125_G2_FS_1_TEMP_P_0_5_0_port, 
      mult_125_G2_FS_1_TEMP_P_0_5_1_port, mult_125_G2_FS_1_TEMP_P_0_5_2_port, 
      mult_125_G2_FS_1_TEMP_P_0_6_0_port, mult_125_G2_FS_1_TEMP_P_0_6_1_port, 
      mult_125_G2_FS_1_TEMP_P_0_6_2_port, mult_125_G2_FS_1_TEMP_P_0_7_0_port, 
      mult_125_G2_FS_1_G_1_0_3_port, mult_125_G2_FS_1_G_1_1_0_port, 
      mult_125_G2_FS_1_G_1_1_1_port, mult_125_G2_FS_1_G_1_1_2_port, 
      mult_125_G2_FS_1_G_2_0_0_port, mult_125_G2_FS_1_TEMP_G_0_3_2_port, 
      mult_125_G2_FS_1_TEMP_G_0_4_1_port, mult_125_G2_FS_1_TEMP_G_0_4_2_port, 
      mult_125_G2_FS_1_TEMP_G_0_5_1_port, mult_125_G2_FS_1_TEMP_G_0_5_2_port, 
      mult_125_G2_FS_1_TEMP_G_0_6_1_port, mult_125_G2_FS_1_TEMP_G_0_6_2_port, 
      mult_125_G2_FS_1_G_n_int_0_3_2_port, mult_125_G2_FS_1_G_n_int_0_3_3_port,
      mult_125_G2_FS_1_G_n_int_0_4_0_port, mult_125_G2_FS_1_G_n_int_0_4_1_port,
      mult_125_G2_FS_1_G_n_int_0_4_2_port, mult_125_G2_FS_1_G_n_int_0_4_3_port,
      mult_125_G2_FS_1_G_n_int_0_5_0_port, mult_125_G2_FS_1_G_n_int_0_5_1_port,
      mult_125_G2_FS_1_G_n_int_0_5_2_port, mult_125_G2_FS_1_G_n_int_0_5_3_port,
      mult_125_G2_FS_1_G_n_int_0_6_0_port, mult_125_G2_FS_1_G_n_int_0_6_1_port,
      mult_125_G2_FS_1_G_n_int_0_6_2_port, mult_125_G2_FS_1_G_n_int_0_6_3_port,
      mult_125_G2_FS_1_G_n_int_0_7_0_port, mult_125_G2_FS_1_G_n_int_0_7_1_port,
      mult_125_G2_FS_1_PG_int_0_3_3_port, mult_125_G2_FS_1_PG_int_0_4_0_port, 
      mult_125_G2_FS_1_PG_int_0_4_1_port, mult_125_G2_FS_1_PG_int_0_4_2_port, 
      mult_125_G2_FS_1_PG_int_0_4_3_port, mult_125_G2_FS_1_PG_int_0_5_0_port, 
      mult_125_G2_FS_1_PG_int_0_5_1_port, mult_125_G2_FS_1_PG_int_0_5_2_port, 
      mult_125_G2_FS_1_PG_int_0_5_3_port, mult_125_G2_FS_1_PG_int_0_6_0_port, 
      mult_125_G2_FS_1_PG_int_0_6_1_port, mult_125_G2_FS_1_PG_int_0_6_2_port, 
      mult_125_G2_FS_1_PG_int_0_6_3_port, mult_125_G2_FS_1_PG_int_0_7_0_port, 
      mult_125_G2_FS_1_PG_int_0_7_1_port, mult_125_G2_A2_14_port, 
      mult_125_G2_A2_15_port, mult_125_G2_A2_16_port, mult_125_G2_A2_17_port, 
      mult_125_G2_A2_18_port, mult_125_G2_A2_19_port, mult_125_G2_A2_20_port, 
      mult_125_G2_A2_21_port, mult_125_G2_A2_22_port, mult_125_G2_A2_23_port, 
      mult_125_G2_A2_24_port, mult_125_G2_A2_25_port, mult_125_G2_A2_26_port, 
      mult_125_G2_A2_27_port, mult_125_G2_A2_28_port, mult_125_G2_A2_29_port, 
      mult_125_G2_A1_0_port, mult_125_G2_A1_1_port, mult_125_G2_A1_2_port, 
      mult_125_G2_A1_3_port, mult_125_G2_A1_4_port, mult_125_G2_A1_5_port, 
      mult_125_G2_A1_6_port, mult_125_G2_A1_7_port, mult_125_G2_A1_8_port, 
      mult_125_G2_A1_9_port, mult_125_G2_A1_10_port, mult_125_G2_A1_11_port, 
      mult_125_G2_A1_12_port, mult_125_G2_A1_13_port, mult_125_G2_A1_14_port, 
      mult_125_G2_A1_15_port, mult_125_G2_A1_16_port, mult_125_G2_A1_17_port, 
      mult_125_G2_A1_18_port, mult_125_G2_A1_19_port, mult_125_G2_A1_20_port, 
      mult_125_G2_A1_21_port, mult_125_G2_A1_22_port, mult_125_G2_A1_23_port, 
      mult_125_G2_A1_24_port, mult_125_G2_A1_25_port, mult_125_G2_A1_26_port, 
      mult_125_G2_A1_27_port, mult_125_G2_A1_28_port, mult_125_G2_A1_29_port, 
      mult_125_G2_ZB, mult_125_G2_ZA, mult_125_G2_QB, mult_125_G2_QA, 
      mult_125_G2_A_notx_0_port, mult_125_G2_A_notx_1_port, 
      mult_125_G2_A_notx_2_port, mult_125_G2_A_notx_3_port, 
      mult_125_G2_A_notx_4_port, mult_125_G2_A_notx_5_port, 
      mult_125_G2_A_notx_6_port, mult_125_G2_A_notx_7_port, 
      mult_125_G2_A_notx_8_port, mult_125_G2_A_notx_9_port, 
      mult_125_G2_A_notx_10_port, mult_125_G2_A_notx_11_port, 
      mult_125_G2_A_notx_12_port, mult_125_G2_A_notx_13_port, 
      mult_125_G2_A_notx_14_port, mult_125_G2_B_notx_0_port, 
      mult_125_G2_B_notx_1_port, mult_125_G2_B_notx_2_port, 
      mult_125_G2_B_notx_3_port, mult_125_G2_B_notx_4_port, 
      mult_125_G2_B_notx_5_port, mult_125_G2_B_notx_6_port, 
      mult_125_G2_B_notx_7_port, mult_125_G2_B_notx_8_port, 
      mult_125_G2_B_notx_9_port, mult_125_G2_B_notx_10_port, 
      mult_125_G2_B_notx_11_port, mult_125_G2_B_notx_12_port, 
      mult_125_G2_B_notx_13_port, mult_125_G2_B_notx_14_port, 
      mult_125_G2_ab_0_1_port, mult_125_G2_ab_0_2_port, mult_125_G2_ab_0_3_port
      , mult_125_G2_ab_0_4_port, mult_125_G2_ab_0_5_port, 
      mult_125_G2_ab_0_6_port, mult_125_G2_ab_0_7_port, mult_125_G2_ab_0_8_port
      , mult_125_G2_ab_0_9_port, mult_125_G2_ab_0_10_port, 
      mult_125_G2_ab_0_11_port, mult_125_G2_ab_0_12_port, 
      mult_125_G2_ab_0_13_port, mult_125_G2_ab_0_14_port, 
      mult_125_G2_ab_0_15_port, mult_125_G2_ab_1_0_port, 
      mult_125_G2_ab_1_1_port, mult_125_G2_ab_1_2_port, mult_125_G2_ab_1_3_port
      , mult_125_G2_ab_1_4_port, mult_125_G2_ab_1_5_port, 
      mult_125_G2_ab_1_6_port, mult_125_G2_ab_1_7_port, mult_125_G2_ab_1_8_port
      , mult_125_G2_ab_1_9_port, mult_125_G2_ab_1_10_port, 
      mult_125_G2_ab_1_11_port, mult_125_G2_ab_1_12_port, 
      mult_125_G2_ab_1_13_port, mult_125_G2_ab_1_14_port, 
      mult_125_G2_ab_1_15_port, mult_125_G2_ab_2_0_port, 
      mult_125_G2_ab_2_1_port, mult_125_G2_ab_2_2_port, mult_125_G2_ab_2_3_port
      , mult_125_G2_ab_2_4_port, mult_125_G2_ab_2_5_port, 
      mult_125_G2_ab_2_6_port, mult_125_G2_ab_2_7_port, mult_125_G2_ab_2_8_port
      , mult_125_G2_ab_2_9_port, mult_125_G2_ab_2_10_port, 
      mult_125_G2_ab_2_11_port, mult_125_G2_ab_2_12_port, 
      mult_125_G2_ab_2_13_port, mult_125_G2_ab_2_14_port, 
      mult_125_G2_ab_2_15_port, mult_125_G2_ab_3_0_port, 
      mult_125_G2_ab_3_1_port, mult_125_G2_ab_3_2_port, mult_125_G2_ab_3_3_port
      , mult_125_G2_ab_3_4_port, mult_125_G2_ab_3_5_port, 
      mult_125_G2_ab_3_6_port, mult_125_G2_ab_3_7_port, mult_125_G2_ab_3_8_port
      , mult_125_G2_ab_3_9_port, mult_125_G2_ab_3_10_port, 
      mult_125_G2_ab_3_11_port, mult_125_G2_ab_3_12_port, 
      mult_125_G2_ab_3_13_port, mult_125_G2_ab_3_14_port, 
      mult_125_G2_ab_3_15_port, mult_125_G2_ab_4_0_port, 
      mult_125_G2_ab_4_1_port, mult_125_G2_ab_4_2_port, mult_125_G2_ab_4_3_port
      , mult_125_G2_ab_4_4_port, mult_125_G2_ab_4_5_port, 
      mult_125_G2_ab_4_6_port, mult_125_G2_ab_4_7_port, mult_125_G2_ab_4_8_port
      , mult_125_G2_ab_4_9_port, mult_125_G2_ab_4_10_port, 
      mult_125_G2_ab_4_11_port, mult_125_G2_ab_4_12_port, 
      mult_125_G2_ab_4_13_port, mult_125_G2_ab_4_14_port, 
      mult_125_G2_ab_4_15_port, mult_125_G2_ab_5_0_port, 
      mult_125_G2_ab_5_1_port, mult_125_G2_ab_5_2_port, mult_125_G2_ab_5_3_port
      , mult_125_G2_ab_5_4_port, mult_125_G2_ab_5_5_port, 
      mult_125_G2_ab_5_6_port, mult_125_G2_ab_5_7_port, mult_125_G2_ab_5_8_port
      , mult_125_G2_ab_5_9_port, mult_125_G2_ab_5_10_port, 
      mult_125_G2_ab_5_11_port, mult_125_G2_ab_5_12_port, 
      mult_125_G2_ab_5_13_port, mult_125_G2_ab_5_14_port, 
      mult_125_G2_ab_5_15_port, mult_125_G2_ab_6_0_port, 
      mult_125_G2_ab_6_1_port, mult_125_G2_ab_6_2_port, mult_125_G2_ab_6_3_port
      , mult_125_G2_ab_6_4_port, mult_125_G2_ab_6_5_port, 
      mult_125_G2_ab_6_6_port, mult_125_G2_ab_6_7_port, mult_125_G2_ab_6_8_port
      , mult_125_G2_ab_6_9_port, mult_125_G2_ab_6_10_port, 
      mult_125_G2_ab_6_11_port, mult_125_G2_ab_6_12_port, 
      mult_125_G2_ab_6_13_port, mult_125_G2_ab_6_14_port, 
      mult_125_G2_ab_6_15_port, mult_125_G2_ab_7_0_port, 
      mult_125_G2_ab_7_1_port, mult_125_G2_ab_7_2_port, mult_125_G2_ab_7_3_port
      , mult_125_G2_ab_7_4_port, mult_125_G2_ab_7_5_port, 
      mult_125_G2_ab_7_6_port, mult_125_G2_ab_7_7_port, mult_125_G2_ab_7_8_port
      , mult_125_G2_ab_7_9_port, mult_125_G2_ab_7_10_port, 
      mult_125_G2_ab_7_11_port, mult_125_G2_ab_7_12_port, 
      mult_125_G2_ab_7_13_port, mult_125_G2_ab_7_14_port, 
      mult_125_G2_ab_7_15_port, mult_125_G2_ab_8_0_port, 
      mult_125_G2_ab_8_1_port, mult_125_G2_ab_8_2_port, mult_125_G2_ab_8_3_port
      , mult_125_G2_ab_8_4_port, mult_125_G2_ab_8_5_port, 
      mult_125_G2_ab_8_6_port, mult_125_G2_ab_8_7_port, mult_125_G2_ab_8_8_port
      , mult_125_G2_ab_8_9_port, mult_125_G2_ab_8_10_port, 
      mult_125_G2_ab_8_11_port, mult_125_G2_ab_8_12_port, 
      mult_125_G2_ab_8_13_port, mult_125_G2_ab_8_14_port, 
      mult_125_G2_ab_8_15_port, mult_125_G2_ab_9_0_port, 
      mult_125_G2_ab_9_1_port, mult_125_G2_ab_9_2_port, mult_125_G2_ab_9_3_port
      , mult_125_G2_ab_9_4_port, mult_125_G2_ab_9_5_port, 
      mult_125_G2_ab_9_6_port, mult_125_G2_ab_9_7_port, mult_125_G2_ab_9_8_port
      , mult_125_G2_ab_9_9_port, mult_125_G2_ab_9_10_port, 
      mult_125_G2_ab_9_11_port, mult_125_G2_ab_9_12_port, 
      mult_125_G2_ab_9_13_port, mult_125_G2_ab_9_14_port, 
      mult_125_G2_ab_9_15_port, mult_125_G2_ab_10_0_port, 
      mult_125_G2_ab_10_1_port, mult_125_G2_ab_10_2_port, 
      mult_125_G2_ab_10_3_port, mult_125_G2_ab_10_4_port, 
      mult_125_G2_ab_10_5_port, mult_125_G2_ab_10_6_port, 
      mult_125_G2_ab_10_7_port, mult_125_G2_ab_10_8_port, 
      mult_125_G2_ab_10_9_port, mult_125_G2_ab_10_10_port, 
      mult_125_G2_ab_10_11_port, mult_125_G2_ab_10_12_port, 
      mult_125_G2_ab_10_13_port, mult_125_G2_ab_10_14_port, 
      mult_125_G2_ab_10_15_port, mult_125_G2_ab_11_0_port, 
      mult_125_G2_ab_11_1_port, mult_125_G2_ab_11_2_port, 
      mult_125_G2_ab_11_3_port, mult_125_G2_ab_11_4_port, 
      mult_125_G2_ab_11_5_port, mult_125_G2_ab_11_6_port, 
      mult_125_G2_ab_11_7_port, mult_125_G2_ab_11_8_port, 
      mult_125_G2_ab_11_9_port, mult_125_G2_ab_11_10_port, 
      mult_125_G2_ab_11_11_port, mult_125_G2_ab_11_12_port, 
      mult_125_G2_ab_11_13_port, mult_125_G2_ab_11_14_port, 
      mult_125_G2_ab_11_15_port, mult_125_G2_ab_12_0_port, 
      mult_125_G2_ab_12_1_port, mult_125_G2_ab_12_2_port, 
      mult_125_G2_ab_12_3_port, mult_125_G2_ab_12_4_port, 
      mult_125_G2_ab_12_5_port, mult_125_G2_ab_12_6_port, 
      mult_125_G2_ab_12_7_port, mult_125_G2_ab_12_8_port, 
      mult_125_G2_ab_12_9_port, mult_125_G2_ab_12_10_port, 
      mult_125_G2_ab_12_11_port, mult_125_G2_ab_12_12_port, 
      mult_125_G2_ab_12_13_port, mult_125_G2_ab_12_14_port, 
      mult_125_G2_ab_12_15_port, mult_125_G2_ab_13_0_port, 
      mult_125_G2_ab_13_1_port, mult_125_G2_ab_13_2_port, 
      mult_125_G2_ab_13_3_port, mult_125_G2_ab_13_4_port, 
      mult_125_G2_ab_13_5_port, mult_125_G2_ab_13_6_port, 
      mult_125_G2_ab_13_7_port, mult_125_G2_ab_13_8_port, 
      mult_125_G2_ab_13_9_port, mult_125_G2_ab_13_10_port, 
      mult_125_G2_ab_13_11_port, mult_125_G2_ab_13_12_port, 
      mult_125_G2_ab_13_13_port, mult_125_G2_ab_13_14_port, 
      mult_125_G2_ab_13_15_port, mult_125_G2_ab_14_0_port, 
      mult_125_G2_ab_14_1_port, mult_125_G2_ab_14_2_port, 
      mult_125_G2_ab_14_3_port, mult_125_G2_ab_14_4_port, 
      mult_125_G2_ab_14_5_port, mult_125_G2_ab_14_6_port, 
      mult_125_G2_ab_14_7_port, mult_125_G2_ab_14_8_port, 
      mult_125_G2_ab_14_9_port, mult_125_G2_ab_14_10_port, 
      mult_125_G2_ab_14_11_port, mult_125_G2_ab_14_12_port, 
      mult_125_G2_ab_14_13_port, mult_125_G2_ab_14_14_port, 
      mult_125_G2_ab_14_15_port, mult_125_G2_ab_15_0_port, 
      mult_125_G2_ab_15_1_port, mult_125_G2_ab_15_2_port, 
      mult_125_G2_ab_15_3_port, mult_125_G2_ab_15_4_port, 
      mult_125_G2_ab_15_5_port, mult_125_G2_ab_15_6_port, 
      mult_125_G2_ab_15_7_port, mult_125_G2_ab_15_8_port, 
      mult_125_G2_ab_15_9_port, mult_125_G2_ab_15_10_port, 
      mult_125_G2_ab_15_11_port, mult_125_G2_ab_15_12_port, 
      mult_125_G2_ab_15_13_port, mult_125_G2_ab_15_14_port, 
      mult_125_G2_ab_15_15_port, mult_125_G2_B_not_0_port, 
      mult_125_G2_B_not_1_port, mult_125_G2_B_not_2_port, 
      mult_125_G2_B_not_3_port, mult_125_G2_B_not_4_port, 
      mult_125_G2_B_not_5_port, mult_125_G2_B_not_6_port, 
      mult_125_G2_B_not_7_port, mult_125_G2_B_not_8_port, 
      mult_125_G2_B_not_9_port, mult_125_G2_B_not_10_port, 
      mult_125_G2_B_not_11_port, mult_125_G2_B_not_12_port, 
      mult_125_G2_B_not_13_port, mult_125_G2_B_not_14_port, 
      mult_125_G2_B_not_15_port, mult_125_G2_A_not_0_port, 
      mult_125_G2_A_not_1_port, mult_125_G2_A_not_2_port, 
      mult_125_G2_A_not_3_port, mult_125_G2_A_not_4_port, 
      mult_125_G2_A_not_5_port, mult_125_G2_A_not_6_port, 
      mult_125_G2_A_not_7_port, mult_125_G2_A_not_8_port, 
      mult_125_G2_A_not_9_port, mult_125_G2_A_not_10_port, 
      mult_125_G2_A_not_11_port, mult_125_G2_A_not_12_port, 
      mult_125_G2_A_not_13_port, mult_125_G2_A_not_14_port, 
      mult_125_G2_A_not_15_port, mult_125_FS_1_C_1_3_3_port, 
      mult_125_FS_1_C_1_4_0_port, mult_125_FS_1_C_1_4_1_port, 
      mult_125_FS_1_C_1_4_2_port, mult_125_FS_1_C_1_4_3_port, 
      mult_125_FS_1_C_1_5_0_port, mult_125_FS_1_C_1_5_1_port, 
      mult_125_FS_1_C_1_5_2_port, mult_125_FS_1_C_1_5_3_port, 
      mult_125_FS_1_C_1_6_0_port, mult_125_FS_1_C_1_6_1_port, 
      mult_125_FS_1_C_1_6_2_port, mult_125_FS_1_C_1_6_3_port, 
      mult_125_FS_1_C_1_7_0_port, mult_125_FS_1_C_1_7_1_port, 
      mult_125_FS_1_P_0_0_1_port, mult_125_FS_1_P_0_0_2_port, 
      mult_125_FS_1_P_0_0_3_port, mult_125_FS_1_P_0_1_1_port, 
      mult_125_FS_1_P_0_1_2_port, mult_125_FS_1_P_0_1_3_port, 
      mult_125_FS_1_P_0_2_1_port, mult_125_FS_1_P_0_2_2_port, 
      mult_125_FS_1_P_0_2_3_port, mult_125_FS_1_P_0_3_1_port, 
      mult_125_FS_1_P_0_3_2_port, mult_125_FS_1_P_0_3_3_port, 
      mult_125_FS_1_P_0_4_1_port, mult_125_FS_1_P_0_4_2_port, 
      mult_125_FS_1_P_0_4_3_port, mult_125_FS_1_P_0_5_1_port, 
      mult_125_FS_1_P_0_5_2_port, mult_125_FS_1_P_0_5_3_port, 
      mult_125_FS_1_P_0_6_1_port, mult_125_FS_1_P_0_6_2_port, 
      mult_125_FS_1_P_0_6_3_port, mult_125_FS_1_P_0_7_1_port, 
      mult_125_FS_1_TEMP_P_0_0_0_port, mult_125_FS_1_TEMP_P_0_1_0_port, 
      mult_125_FS_1_TEMP_P_0_2_0_port, mult_125_FS_1_TEMP_P_0_3_0_port, 
      mult_125_FS_1_TEMP_P_0_4_0_port, mult_125_FS_1_TEMP_P_0_4_1_port, 
      mult_125_FS_1_TEMP_P_0_4_2_port, mult_125_FS_1_TEMP_P_0_5_0_port, 
      mult_125_FS_1_TEMP_P_0_5_1_port, mult_125_FS_1_TEMP_P_0_5_2_port, 
      mult_125_FS_1_TEMP_P_0_6_0_port, mult_125_FS_1_TEMP_P_0_6_1_port, 
      mult_125_FS_1_TEMP_P_0_6_2_port, mult_125_FS_1_TEMP_P_0_7_0_port, 
      mult_125_FS_1_G_1_0_3_port, mult_125_FS_1_G_1_1_0_port, 
      mult_125_FS_1_G_1_1_1_port, mult_125_FS_1_G_1_1_2_port, 
      mult_125_FS_1_G_2_0_0_port, mult_125_FS_1_TEMP_G_0_3_2_port, 
      mult_125_FS_1_TEMP_G_0_4_1_port, mult_125_FS_1_TEMP_G_0_4_2_port, 
      mult_125_FS_1_TEMP_G_0_5_1_port, mult_125_FS_1_TEMP_G_0_5_2_port, 
      mult_125_FS_1_TEMP_G_0_6_1_port, mult_125_FS_1_TEMP_G_0_6_2_port, 
      mult_125_FS_1_G_n_int_0_3_2_port, mult_125_FS_1_G_n_int_0_3_3_port, 
      mult_125_FS_1_G_n_int_0_4_0_port, mult_125_FS_1_G_n_int_0_4_1_port, 
      mult_125_FS_1_G_n_int_0_4_2_port, mult_125_FS_1_G_n_int_0_4_3_port, 
      mult_125_FS_1_G_n_int_0_5_0_port, mult_125_FS_1_G_n_int_0_5_1_port, 
      mult_125_FS_1_G_n_int_0_5_2_port, mult_125_FS_1_G_n_int_0_5_3_port, 
      mult_125_FS_1_G_n_int_0_6_0_port, mult_125_FS_1_G_n_int_0_6_1_port, 
      mult_125_FS_1_G_n_int_0_6_2_port, mult_125_FS_1_G_n_int_0_6_3_port, 
      mult_125_FS_1_G_n_int_0_7_0_port, mult_125_FS_1_G_n_int_0_7_1_port, 
      mult_125_FS_1_PG_int_0_3_3_port, mult_125_FS_1_PG_int_0_4_0_port, 
      mult_125_FS_1_PG_int_0_4_1_port, mult_125_FS_1_PG_int_0_4_2_port, 
      mult_125_FS_1_PG_int_0_4_3_port, mult_125_FS_1_PG_int_0_5_0_port, 
      mult_125_FS_1_PG_int_0_5_1_port, mult_125_FS_1_PG_int_0_5_2_port, 
      mult_125_FS_1_PG_int_0_5_3_port, mult_125_FS_1_PG_int_0_6_0_port, 
      mult_125_FS_1_PG_int_0_6_1_port, mult_125_FS_1_PG_int_0_6_2_port, 
      mult_125_FS_1_PG_int_0_6_3_port, mult_125_FS_1_PG_int_0_7_0_port, 
      mult_125_FS_1_PG_int_0_7_1_port, mult_125_A2_14_port, mult_125_A2_15_port
      , mult_125_A2_16_port, mult_125_A2_17_port, mult_125_A2_18_port, 
      mult_125_A2_19_port, mult_125_A2_20_port, mult_125_A2_21_port, 
      mult_125_A2_22_port, mult_125_A2_23_port, mult_125_A2_24_port, 
      mult_125_A2_25_port, mult_125_A2_26_port, mult_125_A2_27_port, 
      mult_125_A2_28_port, mult_125_A2_29_port, mult_125_A1_0_port, 
      mult_125_A1_1_port, mult_125_A1_2_port, mult_125_A1_3_port, 
      mult_125_A1_4_port, mult_125_A1_5_port, mult_125_A1_6_port, 
      mult_125_A1_7_port, mult_125_A1_8_port, mult_125_A1_9_port, 
      mult_125_A1_10_port, mult_125_A1_11_port, mult_125_A1_12_port, 
      mult_125_A1_13_port, mult_125_A1_14_port, mult_125_A1_15_port, 
      mult_125_A1_16_port, mult_125_A1_17_port, mult_125_A1_18_port, 
      mult_125_A1_19_port, mult_125_A1_20_port, mult_125_A1_21_port, 
      mult_125_A1_22_port, mult_125_A1_23_port, mult_125_A1_24_port, 
      mult_125_A1_25_port, mult_125_A1_26_port, mult_125_A1_27_port, 
      mult_125_A1_28_port, mult_125_A1_29_port, mult_125_ZB, mult_125_ZA, 
      mult_125_QB, mult_125_QA, mult_125_A_notx_0_port, mult_125_A_notx_1_port,
      mult_125_A_notx_2_port, mult_125_A_notx_3_port, mult_125_A_notx_4_port, 
      mult_125_A_notx_5_port, mult_125_A_notx_6_port, mult_125_A_notx_7_port, 
      mult_125_A_notx_8_port, mult_125_A_notx_9_port, mult_125_A_notx_10_port, 
      mult_125_A_notx_11_port, mult_125_A_notx_12_port, mult_125_A_notx_13_port
      , mult_125_A_notx_14_port, mult_125_B_notx_0_port, mult_125_B_notx_1_port
      , mult_125_B_notx_2_port, mult_125_B_notx_3_port, mult_125_B_notx_4_port,
      mult_125_B_notx_5_port, mult_125_B_notx_6_port, mult_125_B_notx_7_port, 
      mult_125_B_notx_8_port, mult_125_B_notx_9_port, mult_125_B_notx_10_port, 
      mult_125_B_notx_11_port, mult_125_B_notx_12_port, mult_125_B_notx_13_port
      , mult_125_B_notx_14_port, mult_125_ab_0_1_port, mult_125_ab_0_2_port, 
      mult_125_ab_0_3_port, mult_125_ab_0_4_port, mult_125_ab_0_5_port, 
      mult_125_ab_0_6_port, mult_125_ab_0_7_port, mult_125_ab_0_8_port, 
      mult_125_ab_0_9_port, mult_125_ab_0_10_port, mult_125_ab_0_11_port, 
      mult_125_ab_0_12_port, mult_125_ab_0_13_port, mult_125_ab_0_14_port, 
      mult_125_ab_0_15_port, mult_125_ab_1_0_port, mult_125_ab_1_1_port, 
      mult_125_ab_1_2_port, mult_125_ab_1_3_port, mult_125_ab_1_4_port, 
      mult_125_ab_1_5_port, mult_125_ab_1_6_port, mult_125_ab_1_7_port, 
      mult_125_ab_1_8_port, mult_125_ab_1_9_port, mult_125_ab_1_10_port, 
      mult_125_ab_1_11_port, mult_125_ab_1_12_port, mult_125_ab_1_13_port, 
      mult_125_ab_1_14_port, mult_125_ab_1_15_port, mult_125_ab_2_0_port, 
      mult_125_ab_2_1_port, mult_125_ab_2_2_port, mult_125_ab_2_3_port, 
      mult_125_ab_2_4_port, mult_125_ab_2_5_port, mult_125_ab_2_6_port, 
      mult_125_ab_2_7_port, mult_125_ab_2_8_port, mult_125_ab_2_9_port, 
      mult_125_ab_2_10_port, mult_125_ab_2_11_port, mult_125_ab_2_12_port, 
      mult_125_ab_2_13_port, mult_125_ab_2_14_port, mult_125_ab_2_15_port, 
      mult_125_ab_3_0_port, mult_125_ab_3_1_port, mult_125_ab_3_2_port, 
      mult_125_ab_3_3_port, mult_125_ab_3_4_port, mult_125_ab_3_5_port, 
      mult_125_ab_3_6_port, mult_125_ab_3_7_port, mult_125_ab_3_8_port, 
      mult_125_ab_3_9_port, mult_125_ab_3_10_port, mult_125_ab_3_11_port, 
      mult_125_ab_3_12_port, mult_125_ab_3_13_port, mult_125_ab_3_14_port, 
      mult_125_ab_3_15_port, mult_125_ab_4_0_port, mult_125_ab_4_1_port, 
      mult_125_ab_4_2_port, mult_125_ab_4_3_port, mult_125_ab_4_4_port, 
      mult_125_ab_4_5_port, mult_125_ab_4_6_port, mult_125_ab_4_7_port, 
      mult_125_ab_4_8_port, mult_125_ab_4_9_port, mult_125_ab_4_10_port, 
      mult_125_ab_4_11_port, mult_125_ab_4_12_port, mult_125_ab_4_13_port, 
      mult_125_ab_4_14_port, mult_125_ab_4_15_port, mult_125_ab_5_0_port, 
      mult_125_ab_5_1_port, mult_125_ab_5_2_port, mult_125_ab_5_3_port, 
      mult_125_ab_5_4_port, mult_125_ab_5_5_port, mult_125_ab_5_6_port, 
      mult_125_ab_5_7_port, mult_125_ab_5_8_port, mult_125_ab_5_9_port, 
      mult_125_ab_5_10_port, mult_125_ab_5_11_port, mult_125_ab_5_12_port, 
      mult_125_ab_5_13_port, mult_125_ab_5_14_port, mult_125_ab_5_15_port, 
      mult_125_ab_6_0_port, mult_125_ab_6_1_port, mult_125_ab_6_2_port, 
      mult_125_ab_6_3_port, mult_125_ab_6_4_port, mult_125_ab_6_5_port, 
      mult_125_ab_6_6_port, mult_125_ab_6_7_port, mult_125_ab_6_8_port, 
      mult_125_ab_6_9_port, mult_125_ab_6_10_port, mult_125_ab_6_11_port, 
      mult_125_ab_6_12_port, mult_125_ab_6_13_port, mult_125_ab_6_14_port, 
      mult_125_ab_6_15_port, mult_125_ab_7_0_port, mult_125_ab_7_1_port, 
      mult_125_ab_7_2_port, mult_125_ab_7_3_port, mult_125_ab_7_4_port, 
      mult_125_ab_7_5_port, mult_125_ab_7_6_port, mult_125_ab_7_7_port, 
      mult_125_ab_7_8_port, mult_125_ab_7_9_port, mult_125_ab_7_10_port, 
      mult_125_ab_7_11_port, mult_125_ab_7_12_port, mult_125_ab_7_13_port, 
      mult_125_ab_7_14_port, mult_125_ab_7_15_port, mult_125_ab_8_0_port, 
      mult_125_ab_8_1_port, mult_125_ab_8_2_port, mult_125_ab_8_3_port, 
      mult_125_ab_8_4_port, mult_125_ab_8_5_port, mult_125_ab_8_6_port, 
      mult_125_ab_8_7_port, mult_125_ab_8_8_port, mult_125_ab_8_9_port, 
      mult_125_ab_8_10_port, mult_125_ab_8_11_port, mult_125_ab_8_12_port, 
      mult_125_ab_8_13_port, mult_125_ab_8_14_port, mult_125_ab_8_15_port, 
      mult_125_ab_9_0_port, mult_125_ab_9_1_port, mult_125_ab_9_2_port, 
      mult_125_ab_9_3_port, mult_125_ab_9_4_port, mult_125_ab_9_5_port, 
      mult_125_ab_9_6_port, mult_125_ab_9_7_port, mult_125_ab_9_8_port, 
      mult_125_ab_9_9_port, mult_125_ab_9_10_port, mult_125_ab_9_11_port, 
      mult_125_ab_9_12_port, mult_125_ab_9_13_port, mult_125_ab_9_14_port, 
      mult_125_ab_9_15_port, mult_125_ab_10_0_port, mult_125_ab_10_1_port, 
      mult_125_ab_10_2_port, mult_125_ab_10_3_port, mult_125_ab_10_4_port, 
      mult_125_ab_10_5_port, mult_125_ab_10_6_port, mult_125_ab_10_7_port, 
      mult_125_ab_10_8_port, mult_125_ab_10_9_port, mult_125_ab_10_10_port, 
      mult_125_ab_10_11_port, mult_125_ab_10_12_port, mult_125_ab_10_13_port, 
      mult_125_ab_10_14_port, mult_125_ab_10_15_port, mult_125_ab_11_0_port, 
      mult_125_ab_11_1_port, mult_125_ab_11_2_port, mult_125_ab_11_3_port, 
      mult_125_ab_11_4_port, mult_125_ab_11_5_port, mult_125_ab_11_6_port, 
      mult_125_ab_11_7_port, mult_125_ab_11_8_port, mult_125_ab_11_9_port, 
      mult_125_ab_11_10_port, mult_125_ab_11_11_port, mult_125_ab_11_12_port, 
      mult_125_ab_11_13_port, mult_125_ab_11_14_port, mult_125_ab_11_15_port, 
      mult_125_ab_12_0_port, mult_125_ab_12_1_port, mult_125_ab_12_2_port, 
      mult_125_ab_12_3_port, mult_125_ab_12_4_port, mult_125_ab_12_5_port, 
      mult_125_ab_12_6_port, mult_125_ab_12_7_port, mult_125_ab_12_8_port, 
      mult_125_ab_12_9_port, mult_125_ab_12_10_port, mult_125_ab_12_11_port, 
      mult_125_ab_12_12_port, mult_125_ab_12_13_port, mult_125_ab_12_14_port, 
      mult_125_ab_12_15_port, mult_125_ab_13_0_port, mult_125_ab_13_1_port, 
      mult_125_ab_13_2_port, mult_125_ab_13_3_port, mult_125_ab_13_4_port, 
      mult_125_ab_13_5_port, mult_125_ab_13_6_port, mult_125_ab_13_7_port, 
      mult_125_ab_13_8_port, mult_125_ab_13_9_port, mult_125_ab_13_10_port, 
      mult_125_ab_13_11_port, mult_125_ab_13_12_port, mult_125_ab_13_13_port, 
      mult_125_ab_13_14_port, mult_125_ab_13_15_port, mult_125_ab_14_0_port, 
      mult_125_ab_14_1_port, mult_125_ab_14_2_port, mult_125_ab_14_3_port, 
      mult_125_ab_14_4_port, mult_125_ab_14_5_port, mult_125_ab_14_6_port, 
      mult_125_ab_14_7_port, mult_125_ab_14_8_port, mult_125_ab_14_9_port, 
      mult_125_ab_14_10_port, mult_125_ab_14_11_port, mult_125_ab_14_12_port, 
      mult_125_ab_14_13_port, mult_125_ab_14_14_port, mult_125_ab_14_15_port, 
      mult_125_ab_15_0_port, mult_125_ab_15_1_port, mult_125_ab_15_2_port, 
      mult_125_ab_15_3_port, mult_125_ab_15_4_port, mult_125_ab_15_5_port, 
      mult_125_ab_15_6_port, mult_125_ab_15_7_port, mult_125_ab_15_8_port, 
      mult_125_ab_15_9_port, mult_125_ab_15_10_port, mult_125_ab_15_11_port, 
      mult_125_ab_15_12_port, mult_125_ab_15_13_port, mult_125_ab_15_14_port, 
      mult_125_ab_15_15_port, mult_125_B_not_0_port, mult_125_B_not_1_port, 
      mult_125_B_not_2_port, mult_125_B_not_3_port, mult_125_B_not_4_port, 
      mult_125_B_not_5_port, mult_125_B_not_6_port, mult_125_B_not_7_port, 
      mult_125_B_not_8_port, mult_125_B_not_9_port, mult_125_B_not_10_port, 
      mult_125_B_not_11_port, mult_125_B_not_12_port, mult_125_B_not_13_port, 
      mult_125_B_not_14_port, mult_125_B_not_15_port, mult_125_A_not_0_port, 
      mult_125_A_not_1_port, mult_125_A_not_2_port, mult_125_A_not_3_port, 
      mult_125_A_not_4_port, mult_125_A_not_5_port, mult_125_A_not_6_port, 
      mult_125_A_not_7_port, mult_125_A_not_8_port, mult_125_A_not_9_port, 
      mult_125_A_not_10_port, mult_125_A_not_11_port, mult_125_A_not_12_port, 
      mult_125_A_not_13_port, mult_125_A_not_14_port, mult_125_A_not_15_port, 
      mult_125_G4_FS_1_C_1_3_3_port, mult_125_G4_FS_1_C_1_4_0_port, 
      mult_125_G4_FS_1_C_1_4_1_port, mult_125_G4_FS_1_C_1_4_2_port, 
      mult_125_G4_FS_1_C_1_4_3_port, mult_125_G4_FS_1_C_1_5_0_port, 
      mult_125_G4_FS_1_C_1_5_1_port, mult_125_G4_FS_1_C_1_5_2_port, 
      mult_125_G4_FS_1_C_1_5_3_port, mult_125_G4_FS_1_C_1_6_0_port, 
      mult_125_G4_FS_1_C_1_6_1_port, mult_125_G4_FS_1_C_1_6_2_port, 
      mult_125_G4_FS_1_C_1_6_3_port, mult_125_G4_FS_1_C_1_7_0_port, 
      mult_125_G4_FS_1_C_1_7_1_port, mult_125_G4_FS_1_P_0_0_1_port, 
      mult_125_G4_FS_1_P_0_0_2_port, mult_125_G4_FS_1_P_0_0_3_port, 
      mult_125_G4_FS_1_P_0_1_1_port, mult_125_G4_FS_1_P_0_1_2_port, 
      mult_125_G4_FS_1_P_0_1_3_port, mult_125_G4_FS_1_P_0_2_1_port, 
      mult_125_G4_FS_1_P_0_2_2_port, mult_125_G4_FS_1_P_0_2_3_port, 
      mult_125_G4_FS_1_P_0_3_1_port, mult_125_G4_FS_1_P_0_3_2_port, 
      mult_125_G4_FS_1_P_0_3_3_port, mult_125_G4_FS_1_P_0_4_1_port, 
      mult_125_G4_FS_1_P_0_4_2_port, mult_125_G4_FS_1_P_0_4_3_port, 
      mult_125_G4_FS_1_P_0_5_1_port, mult_125_G4_FS_1_P_0_5_2_port, 
      mult_125_G4_FS_1_P_0_5_3_port, mult_125_G4_FS_1_P_0_6_1_port, 
      mult_125_G4_FS_1_P_0_6_2_port, mult_125_G4_FS_1_P_0_6_3_port, 
      mult_125_G4_FS_1_P_0_7_1_port, mult_125_G4_FS_1_TEMP_P_0_0_0_port, 
      mult_125_G4_FS_1_TEMP_P_0_1_0_port, mult_125_G4_FS_1_TEMP_P_0_2_0_port, 
      mult_125_G4_FS_1_TEMP_P_0_3_0_port, mult_125_G4_FS_1_TEMP_P_0_4_0_port, 
      mult_125_G4_FS_1_TEMP_P_0_4_1_port, mult_125_G4_FS_1_TEMP_P_0_4_2_port, 
      mult_125_G4_FS_1_TEMP_P_0_5_0_port, mult_125_G4_FS_1_TEMP_P_0_5_1_port, 
      mult_125_G4_FS_1_TEMP_P_0_5_2_port, mult_125_G4_FS_1_TEMP_P_0_6_0_port, 
      mult_125_G4_FS_1_TEMP_P_0_6_1_port, mult_125_G4_FS_1_TEMP_P_0_6_2_port, 
      mult_125_G4_FS_1_TEMP_P_0_7_0_port, mult_125_G4_FS_1_G_1_0_3_port, 
      mult_125_G4_FS_1_G_1_1_0_port, mult_125_G4_FS_1_G_1_1_1_port, 
      mult_125_G4_FS_1_G_1_1_2_port, mult_125_G4_FS_1_G_2_0_0_port, 
      mult_125_G4_FS_1_TEMP_G_0_3_2_port, mult_125_G4_FS_1_TEMP_G_0_4_1_port, 
      mult_125_G4_FS_1_TEMP_G_0_4_2_port, mult_125_G4_FS_1_TEMP_G_0_5_1_port, 
      mult_125_G4_FS_1_TEMP_G_0_5_2_port, mult_125_G4_FS_1_TEMP_G_0_6_1_port, 
      mult_125_G4_FS_1_TEMP_G_0_6_2_port, mult_125_G4_FS_1_G_n_int_0_3_2_port, 
      mult_125_G4_FS_1_G_n_int_0_3_3_port, mult_125_G4_FS_1_G_n_int_0_4_0_port,
      mult_125_G4_FS_1_G_n_int_0_4_1_port, mult_125_G4_FS_1_G_n_int_0_4_2_port,
      mult_125_G4_FS_1_G_n_int_0_4_3_port, mult_125_G4_FS_1_G_n_int_0_5_0_port,
      mult_125_G4_FS_1_G_n_int_0_5_1_port, mult_125_G4_FS_1_G_n_int_0_5_2_port,
      mult_125_G4_FS_1_G_n_int_0_5_3_port, mult_125_G4_FS_1_G_n_int_0_6_0_port,
      mult_125_G4_FS_1_G_n_int_0_6_1_port, mult_125_G4_FS_1_G_n_int_0_6_2_port,
      mult_125_G4_FS_1_G_n_int_0_6_3_port, mult_125_G4_FS_1_G_n_int_0_7_0_port,
      mult_125_G4_FS_1_G_n_int_0_7_1_port, mult_125_G4_FS_1_PG_int_0_3_3_port, 
      mult_125_G4_FS_1_PG_int_0_4_0_port, mult_125_G4_FS_1_PG_int_0_4_1_port, 
      mult_125_G4_FS_1_PG_int_0_4_2_port, mult_125_G4_FS_1_PG_int_0_4_3_port, 
      mult_125_G4_FS_1_PG_int_0_5_0_port, mult_125_G4_FS_1_PG_int_0_5_1_port, 
      mult_125_G4_FS_1_PG_int_0_5_2_port, mult_125_G4_FS_1_PG_int_0_5_3_port, 
      mult_125_G4_FS_1_PG_int_0_6_0_port, mult_125_G4_FS_1_PG_int_0_6_1_port, 
      mult_125_G4_FS_1_PG_int_0_6_2_port, mult_125_G4_FS_1_PG_int_0_6_3_port, 
      mult_125_G4_FS_1_PG_int_0_7_0_port, mult_125_G4_FS_1_PG_int_0_7_1_port, 
      mult_125_G4_A2_14_port, mult_125_G4_A2_15_port, mult_125_G4_A2_16_port, 
      mult_125_G4_A2_17_port, mult_125_G4_A2_18_port, mult_125_G4_A2_19_port, 
      mult_125_G4_A2_20_port, mult_125_G4_A2_21_port, mult_125_G4_A2_22_port, 
      mult_125_G4_A2_23_port, mult_125_G4_A2_24_port, mult_125_G4_A2_25_port, 
      mult_125_G4_A2_26_port, mult_125_G4_A2_27_port, mult_125_G4_A2_28_port, 
      mult_125_G4_A2_29_port, mult_125_G4_A1_0_port, mult_125_G4_A1_1_port, 
      mult_125_G4_A1_2_port, mult_125_G4_A1_3_port, mult_125_G4_A1_4_port, 
      mult_125_G4_A1_5_port, mult_125_G4_A1_6_port, mult_125_G4_A1_7_port, 
      mult_125_G4_A1_8_port, mult_125_G4_A1_9_port, mult_125_G4_A1_10_port, 
      mult_125_G4_A1_11_port, mult_125_G4_A1_12_port, mult_125_G4_A1_13_port, 
      mult_125_G4_A1_14_port, mult_125_G4_A1_15_port, mult_125_G4_A1_16_port, 
      mult_125_G4_A1_17_port, mult_125_G4_A1_18_port, mult_125_G4_A1_19_port, 
      mult_125_G4_A1_20_port, mult_125_G4_A1_21_port, mult_125_G4_A1_22_port, 
      mult_125_G4_A1_23_port, mult_125_G4_A1_24_port, mult_125_G4_A1_25_port, 
      mult_125_G4_A1_26_port, mult_125_G4_A1_27_port, mult_125_G4_A1_28_port, 
      mult_125_G4_A1_29_port, mult_125_G4_ZB, mult_125_G4_ZA, mult_125_G4_QB, 
      mult_125_G4_QA, mult_125_G4_A_notx_0_port, mult_125_G4_A_notx_1_port, 
      mult_125_G4_A_notx_2_port, mult_125_G4_A_notx_3_port, 
      mult_125_G4_A_notx_4_port, mult_125_G4_A_notx_5_port, 
      mult_125_G4_A_notx_6_port, mult_125_G4_A_notx_7_port, 
      mult_125_G4_A_notx_8_port, mult_125_G4_A_notx_9_port, 
      mult_125_G4_A_notx_10_port, mult_125_G4_A_notx_11_port, 
      mult_125_G4_A_notx_12_port, mult_125_G4_A_notx_13_port, 
      mult_125_G4_A_notx_14_port, mult_125_G4_B_notx_0_port, 
      mult_125_G4_B_notx_1_port, mult_125_G4_B_notx_2_port, 
      mult_125_G4_B_notx_3_port, mult_125_G4_B_notx_4_port, 
      mult_125_G4_B_notx_5_port, mult_125_G4_B_notx_6_port, 
      mult_125_G4_B_notx_7_port, mult_125_G4_B_notx_8_port, 
      mult_125_G4_B_notx_9_port, mult_125_G4_B_notx_10_port, 
      mult_125_G4_B_notx_11_port, mult_125_G4_B_notx_12_port, 
      mult_125_G4_B_notx_13_port, mult_125_G4_B_notx_14_port, 
      mult_125_G4_ab_0_1_port, mult_125_G4_ab_0_2_port, mult_125_G4_ab_0_3_port
      , mult_125_G4_ab_0_4_port, mult_125_G4_ab_0_5_port, 
      mult_125_G4_ab_0_6_port, mult_125_G4_ab_0_7_port, mult_125_G4_ab_0_8_port
      , mult_125_G4_ab_0_9_port, mult_125_G4_ab_0_10_port, 
      mult_125_G4_ab_0_11_port, mult_125_G4_ab_0_12_port, 
      mult_125_G4_ab_0_13_port, mult_125_G4_ab_0_14_port, 
      mult_125_G4_ab_0_15_port, mult_125_G4_ab_1_0_port, 
      mult_125_G4_ab_1_1_port, mult_125_G4_ab_1_2_port, mult_125_G4_ab_1_3_port
      , mult_125_G4_ab_1_4_port, mult_125_G4_ab_1_5_port, 
      mult_125_G4_ab_1_6_port, mult_125_G4_ab_1_7_port, mult_125_G4_ab_1_8_port
      , mult_125_G4_ab_1_9_port, mult_125_G4_ab_1_10_port, 
      mult_125_G4_ab_1_11_port, mult_125_G4_ab_1_12_port, 
      mult_125_G4_ab_1_13_port, mult_125_G4_ab_1_14_port, 
      mult_125_G4_ab_1_15_port, mult_125_G4_ab_2_0_port, 
      mult_125_G4_ab_2_1_port, mult_125_G4_ab_2_2_port, mult_125_G4_ab_2_3_port
      , mult_125_G4_ab_2_4_port, mult_125_G4_ab_2_5_port, 
      mult_125_G4_ab_2_6_port, mult_125_G4_ab_2_7_port, mult_125_G4_ab_2_8_port
      , mult_125_G4_ab_2_9_port, mult_125_G4_ab_2_10_port, 
      mult_125_G4_ab_2_11_port, mult_125_G4_ab_2_12_port, 
      mult_125_G4_ab_2_13_port, mult_125_G4_ab_2_14_port, 
      mult_125_G4_ab_2_15_port, mult_125_G4_ab_3_0_port, 
      mult_125_G4_ab_3_1_port, mult_125_G4_ab_3_2_port, mult_125_G4_ab_3_3_port
      , mult_125_G4_ab_3_4_port, mult_125_G4_ab_3_5_port, 
      mult_125_G4_ab_3_6_port, mult_125_G4_ab_3_7_port, mult_125_G4_ab_3_8_port
      , mult_125_G4_ab_3_9_port, mult_125_G4_ab_3_10_port, 
      mult_125_G4_ab_3_11_port, mult_125_G4_ab_3_12_port, 
      mult_125_G4_ab_3_13_port, mult_125_G4_ab_3_14_port, 
      mult_125_G4_ab_3_15_port, mult_125_G4_ab_4_0_port, 
      mult_125_G4_ab_4_1_port, mult_125_G4_ab_4_2_port, mult_125_G4_ab_4_3_port
      , mult_125_G4_ab_4_4_port, mult_125_G4_ab_4_5_port, 
      mult_125_G4_ab_4_6_port, mult_125_G4_ab_4_7_port, mult_125_G4_ab_4_8_port
      , mult_125_G4_ab_4_9_port, mult_125_G4_ab_4_10_port, 
      mult_125_G4_ab_4_11_port, mult_125_G4_ab_4_12_port, 
      mult_125_G4_ab_4_13_port, mult_125_G4_ab_4_14_port, 
      mult_125_G4_ab_4_15_port, mult_125_G4_ab_5_0_port, 
      mult_125_G4_ab_5_1_port, mult_125_G4_ab_5_2_port, mult_125_G4_ab_5_3_port
      , mult_125_G4_ab_5_4_port, mult_125_G4_ab_5_5_port, 
      mult_125_G4_ab_5_6_port, mult_125_G4_ab_5_7_port, mult_125_G4_ab_5_8_port
      , mult_125_G4_ab_5_9_port, mult_125_G4_ab_5_10_port, 
      mult_125_G4_ab_5_11_port, mult_125_G4_ab_5_12_port, 
      mult_125_G4_ab_5_13_port, mult_125_G4_ab_5_14_port, 
      mult_125_G4_ab_5_15_port, mult_125_G4_ab_6_0_port, 
      mult_125_G4_ab_6_1_port, mult_125_G4_ab_6_2_port, mult_125_G4_ab_6_3_port
      , mult_125_G4_ab_6_4_port, mult_125_G4_ab_6_5_port, 
      mult_125_G4_ab_6_6_port, mult_125_G4_ab_6_7_port, mult_125_G4_ab_6_8_port
      , mult_125_G4_ab_6_9_port, mult_125_G4_ab_6_10_port, 
      mult_125_G4_ab_6_11_port, mult_125_G4_ab_6_12_port, 
      mult_125_G4_ab_6_13_port, mult_125_G4_ab_6_14_port, 
      mult_125_G4_ab_6_15_port, mult_125_G4_ab_7_0_port, 
      mult_125_G4_ab_7_1_port, mult_125_G4_ab_7_2_port, mult_125_G4_ab_7_3_port
      , mult_125_G4_ab_7_4_port, mult_125_G4_ab_7_5_port, 
      mult_125_G4_ab_7_6_port, mult_125_G4_ab_7_7_port, mult_125_G4_ab_7_8_port
      , mult_125_G4_ab_7_9_port, mult_125_G4_ab_7_10_port, 
      mult_125_G4_ab_7_11_port, mult_125_G4_ab_7_12_port, 
      mult_125_G4_ab_7_13_port, mult_125_G4_ab_7_14_port, 
      mult_125_G4_ab_7_15_port, mult_125_G4_ab_8_0_port, 
      mult_125_G4_ab_8_1_port, mult_125_G4_ab_8_2_port, mult_125_G4_ab_8_3_port
      , mult_125_G4_ab_8_4_port, mult_125_G4_ab_8_5_port, 
      mult_125_G4_ab_8_6_port, mult_125_G4_ab_8_7_port, mult_125_G4_ab_8_8_port
      , mult_125_G4_ab_8_9_port, mult_125_G4_ab_8_10_port, 
      mult_125_G4_ab_8_11_port, mult_125_G4_ab_8_12_port, 
      mult_125_G4_ab_8_13_port, mult_125_G4_ab_8_14_port, 
      mult_125_G4_ab_8_15_port, mult_125_G4_ab_9_0_port, 
      mult_125_G4_ab_9_1_port, mult_125_G4_ab_9_2_port, mult_125_G4_ab_9_3_port
      , mult_125_G4_ab_9_4_port, mult_125_G4_ab_9_5_port, 
      mult_125_G4_ab_9_6_port, mult_125_G4_ab_9_7_port, mult_125_G4_ab_9_8_port
      , mult_125_G4_ab_9_9_port, mult_125_G4_ab_9_10_port, 
      mult_125_G4_ab_9_11_port, mult_125_G4_ab_9_12_port, 
      mult_125_G4_ab_9_13_port, mult_125_G4_ab_9_14_port, 
      mult_125_G4_ab_9_15_port, mult_125_G4_ab_10_0_port, 
      mult_125_G4_ab_10_1_port, mult_125_G4_ab_10_2_port, 
      mult_125_G4_ab_10_3_port, mult_125_G4_ab_10_4_port, 
      mult_125_G4_ab_10_5_port, mult_125_G4_ab_10_6_port, 
      mult_125_G4_ab_10_7_port, mult_125_G4_ab_10_8_port, 
      mult_125_G4_ab_10_9_port, mult_125_G4_ab_10_10_port, 
      mult_125_G4_ab_10_11_port, mult_125_G4_ab_10_12_port, 
      mult_125_G4_ab_10_13_port, mult_125_G4_ab_10_14_port, 
      mult_125_G4_ab_10_15_port, mult_125_G4_ab_11_0_port, 
      mult_125_G4_ab_11_1_port, mult_125_G4_ab_11_2_port, 
      mult_125_G4_ab_11_3_port, mult_125_G4_ab_11_4_port, 
      mult_125_G4_ab_11_5_port, mult_125_G4_ab_11_6_port, 
      mult_125_G4_ab_11_7_port, mult_125_G4_ab_11_8_port, 
      mult_125_G4_ab_11_9_port, mult_125_G4_ab_11_10_port, 
      mult_125_G4_ab_11_11_port, mult_125_G4_ab_11_12_port, 
      mult_125_G4_ab_11_13_port, mult_125_G4_ab_11_14_port, 
      mult_125_G4_ab_11_15_port, mult_125_G4_ab_12_0_port, 
      mult_125_G4_ab_12_1_port, mult_125_G4_ab_12_2_port, 
      mult_125_G4_ab_12_3_port, mult_125_G4_ab_12_4_port, 
      mult_125_G4_ab_12_5_port, mult_125_G4_ab_12_6_port, 
      mult_125_G4_ab_12_7_port, mult_125_G4_ab_12_8_port, 
      mult_125_G4_ab_12_9_port, mult_125_G4_ab_12_10_port, 
      mult_125_G4_ab_12_11_port, mult_125_G4_ab_12_12_port, 
      mult_125_G4_ab_12_13_port, mult_125_G4_ab_12_14_port, 
      mult_125_G4_ab_12_15_port, mult_125_G4_ab_13_0_port, 
      mult_125_G4_ab_13_1_port, mult_125_G4_ab_13_2_port, 
      mult_125_G4_ab_13_3_port, mult_125_G4_ab_13_4_port, 
      mult_125_G4_ab_13_5_port, mult_125_G4_ab_13_6_port, 
      mult_125_G4_ab_13_7_port, mult_125_G4_ab_13_8_port, 
      mult_125_G4_ab_13_9_port, mult_125_G4_ab_13_10_port, 
      mult_125_G4_ab_13_11_port, mult_125_G4_ab_13_12_port, 
      mult_125_G4_ab_13_13_port, mult_125_G4_ab_13_14_port, 
      mult_125_G4_ab_13_15_port, mult_125_G4_ab_14_0_port, 
      mult_125_G4_ab_14_1_port, mult_125_G4_ab_14_2_port, 
      mult_125_G4_ab_14_3_port, mult_125_G4_ab_14_4_port, 
      mult_125_G4_ab_14_5_port, mult_125_G4_ab_14_6_port, 
      mult_125_G4_ab_14_7_port, mult_125_G4_ab_14_8_port, 
      mult_125_G4_ab_14_9_port, mult_125_G4_ab_14_10_port, 
      mult_125_G4_ab_14_11_port, mult_125_G4_ab_14_12_port, 
      mult_125_G4_ab_14_13_port, mult_125_G4_ab_14_14_port, 
      mult_125_G4_ab_14_15_port, mult_125_G4_ab_15_0_port, 
      mult_125_G4_ab_15_1_port, mult_125_G4_ab_15_2_port, 
      mult_125_G4_ab_15_3_port, mult_125_G4_ab_15_4_port, 
      mult_125_G4_ab_15_5_port, mult_125_G4_ab_15_6_port, 
      mult_125_G4_ab_15_7_port, mult_125_G4_ab_15_8_port, 
      mult_125_G4_ab_15_9_port, mult_125_G4_ab_15_10_port, 
      mult_125_G4_ab_15_11_port, mult_125_G4_ab_15_12_port, 
      mult_125_G4_ab_15_13_port, mult_125_G4_ab_15_14_port, 
      mult_125_G4_ab_15_15_port, mult_125_G4_B_not_0_port, 
      mult_125_G4_B_not_1_port, mult_125_G4_B_not_2_port, 
      mult_125_G4_B_not_3_port, mult_125_G4_B_not_4_port, 
      mult_125_G4_B_not_5_port, mult_125_G4_B_not_6_port, 
      mult_125_G4_B_not_7_port, mult_125_G4_B_not_8_port, 
      mult_125_G4_B_not_9_port, mult_125_G4_B_not_10_port, 
      mult_125_G4_B_not_11_port, mult_125_G4_B_not_12_port, 
      mult_125_G4_B_not_13_port, mult_125_G4_B_not_14_port, 
      mult_125_G4_B_not_15_port, mult_125_G4_A_not_0_port, 
      mult_125_G4_A_not_1_port, mult_125_G4_A_not_2_port, 
      mult_125_G4_A_not_3_port, mult_125_G4_A_not_4_port, 
      mult_125_G4_A_not_5_port, mult_125_G4_A_not_6_port, 
      mult_125_G4_A_not_7_port, mult_125_G4_A_not_8_port, 
      mult_125_G4_A_not_9_port, mult_125_G4_A_not_10_port, 
      mult_125_G4_A_not_11_port, mult_125_G4_A_not_12_port, 
      mult_125_G4_A_not_13_port, mult_125_G4_A_not_14_port, 
      mult_125_G4_A_not_15_port, n240, n241, n242, n243, n244, n245, n246, n247
      , n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
      n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, 
      n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
      n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
      n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
      n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
      n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
      n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, 
      n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, 
      n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
      n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, 
      n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, 
      n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
      n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
      n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, 
      n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, 
      n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, 
      n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, 
      n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, 
      n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, 
      n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
      n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
      n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
      n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
      n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, 
      n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, 
      n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
      n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, 
      n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, 
      n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, 
      n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
      n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, 
      n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, 
      n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, 
      n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, 
      n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, 
      n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, 
      n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, 
      n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, 
      n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, 
      n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, 
      n6033, n6034, n6035 : std_logic;

begin
   ready_x_out <= ready_x_out_port;
   ready_h_out <= ready_h_out_port;
   valid_out <= valid_out_port;
   
   adder_mem_array_reg_3_0_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_0_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_0_port);
   adder_mem_array_reg_3_1_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_1_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_1_port);
   adder_mem_array_reg_3_2_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_2_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_2_port);
   adder_mem_array_reg_3_3_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_3_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_3_port);
   adder_mem_array_reg_3_4_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_4_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_4_port);
   adder_mem_array_reg_3_5_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_5_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_5_port);
   adder_mem_array_reg_3_6_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_6_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_6_port);
   adder_mem_array_reg_3_7_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_7_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_7_port);
   adder_mem_array_reg_3_8_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_8_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_8_port);
   adder_mem_array_reg_3_9_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_9_port, gclk => clk, asyncrsthl =>
                           rst, q => adder_mem_array_3_9_port);
   adder_mem_array_reg_3_10_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_10_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_10_port);
   adder_mem_array_reg_3_11_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_11_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_11_port);
   adder_mem_array_reg_3_12_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_12_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_12_port);
   adder_mem_array_reg_3_13_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_13_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_13_port);
   adder_mem_array_reg_3_14_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_14_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_14_port);
   adder_mem_array_reg_3_15_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_15_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_15_port);
   adder_mem_array_reg_3_16_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_16_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_16_port);
   adder_mem_array_reg_3_17_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_17_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_17_port);
   adder_mem_array_reg_3_18_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_18_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_18_port);
   adder_mem_array_reg_3_19_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_19_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_19_port);
   adder_mem_array_reg_3_20_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_20_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_20_port);
   adder_mem_array_reg_3_21_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_21_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_21_port);
   adder_mem_array_reg_3_22_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_22_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_22_port);
   adder_mem_array_reg_3_23_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_23_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_23_port);
   adder_mem_array_reg_3_24_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_24_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_24_port);
   adder_mem_array_reg_3_25_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_25_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_25_port);
   adder_mem_array_reg_3_26_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_26_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_26_port);
   adder_mem_array_reg_3_27_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_27_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_27_port);
   adder_mem_array_reg_3_28_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_28_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_28_port);
   adder_mem_array_reg_3_29_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_29_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_29_port);
   adder_mem_array_reg_3_30_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_30_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_30_port);
   adder_mem_array_reg_3_32_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_31_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_32_port);
   adder_mem_array_reg_3_31_inst : dff_asyncrsthl port map( d => 
                           multiplier_sigs_3_31_port, gclk => clk, asyncrsthl 
                           => rst, q => adder_mem_array_3_31_port);
   adder_mem_array_reg_2_0_inst : dff_asyncrsthl port map( d => N72, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_0_port);
   adder_mem_array_reg_2_1_inst : dff_asyncrsthl port map( d => N73, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_1_port);
   adder_mem_array_reg_2_2_inst : dff_asyncrsthl port map( d => N74, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_2_port);
   adder_mem_array_reg_2_3_inst : dff_asyncrsthl port map( d => N75, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_3_port);
   adder_mem_array_reg_2_4_inst : dff_asyncrsthl port map( d => N76, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_4_port);
   adder_mem_array_reg_2_5_inst : dff_asyncrsthl port map( d => N77, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_5_port);
   adder_mem_array_reg_2_6_inst : dff_asyncrsthl port map( d => N78, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_6_port);
   adder_mem_array_reg_2_7_inst : dff_asyncrsthl port map( d => N79, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_7_port);
   adder_mem_array_reg_2_8_inst : dff_asyncrsthl port map( d => N80, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_8_port);
   adder_mem_array_reg_2_9_inst : dff_asyncrsthl port map( d => N81, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_9_port);
   adder_mem_array_reg_2_10_inst : dff_asyncrsthl port map( d => N82, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_10_port);
   adder_mem_array_reg_2_11_inst : dff_asyncrsthl port map( d => N83, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_11_port);
   adder_mem_array_reg_2_12_inst : dff_asyncrsthl port map( d => N84, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_12_port);
   adder_mem_array_reg_2_13_inst : dff_asyncrsthl port map( d => N85, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_13_port);
   adder_mem_array_reg_2_14_inst : dff_asyncrsthl port map( d => N86, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_14_port);
   adder_mem_array_reg_2_15_inst : dff_asyncrsthl port map( d => N87, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_15_port);
   adder_mem_array_reg_2_16_inst : dff_asyncrsthl port map( d => N88, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_16_port);
   adder_mem_array_reg_2_17_inst : dff_asyncrsthl port map( d => N89, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_17_port);
   adder_mem_array_reg_2_18_inst : dff_asyncrsthl port map( d => N90, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_18_port);
   adder_mem_array_reg_2_19_inst : dff_asyncrsthl port map( d => N91, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_19_port);
   adder_mem_array_reg_2_20_inst : dff_asyncrsthl port map( d => N92, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_20_port);
   adder_mem_array_reg_2_21_inst : dff_asyncrsthl port map( d => N93, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_21_port);
   adder_mem_array_reg_2_22_inst : dff_asyncrsthl port map( d => N94, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_22_port);
   adder_mem_array_reg_2_23_inst : dff_asyncrsthl port map( d => N95, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_23_port);
   adder_mem_array_reg_2_24_inst : dff_asyncrsthl port map( d => N96, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_24_port);
   adder_mem_array_reg_2_25_inst : dff_asyncrsthl port map( d => N97, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_25_port);
   adder_mem_array_reg_2_26_inst : dff_asyncrsthl port map( d => N98, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_26_port);
   adder_mem_array_reg_2_27_inst : dff_asyncrsthl port map( d => N99, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_27_port);
   adder_mem_array_reg_2_28_inst : dff_asyncrsthl port map( d => N100, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_28_port);
   adder_mem_array_reg_2_29_inst : dff_asyncrsthl port map( d => N101, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_29_port);
   adder_mem_array_reg_2_30_inst : dff_asyncrsthl port map( d => N102, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_30_port);
   adder_mem_array_reg_2_31_inst : dff_asyncrsthl port map( d => N103, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_31_port);
   adder_mem_array_reg_2_32_inst : dff_asyncrsthl port map( d => N104, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_2_32_port);
   adder_mem_array_reg_1_0_inst : dff_asyncrsthl port map( d => N39, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_0_port);
   adder_mem_array_reg_1_1_inst : dff_asyncrsthl port map( d => N40, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_1_port);
   adder_mem_array_reg_1_2_inst : dff_asyncrsthl port map( d => N41, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_2_port);
   adder_mem_array_reg_1_3_inst : dff_asyncrsthl port map( d => N42, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_3_port);
   adder_mem_array_reg_1_4_inst : dff_asyncrsthl port map( d => N43, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_4_port);
   adder_mem_array_reg_1_5_inst : dff_asyncrsthl port map( d => N44, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_5_port);
   adder_mem_array_reg_1_6_inst : dff_asyncrsthl port map( d => N45, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_6_port);
   adder_mem_array_reg_1_7_inst : dff_asyncrsthl port map( d => N46, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_7_port);
   adder_mem_array_reg_1_8_inst : dff_asyncrsthl port map( d => N47, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_8_port);
   adder_mem_array_reg_1_9_inst : dff_asyncrsthl port map( d => N48, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_9_port);
   adder_mem_array_reg_1_10_inst : dff_asyncrsthl port map( d => N49, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_10_port);
   adder_mem_array_reg_1_11_inst : dff_asyncrsthl port map( d => N50, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_11_port);
   adder_mem_array_reg_1_12_inst : dff_asyncrsthl port map( d => N51, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_12_port);
   adder_mem_array_reg_1_13_inst : dff_asyncrsthl port map( d => N52, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_13_port);
   adder_mem_array_reg_1_14_inst : dff_asyncrsthl port map( d => N53, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_14_port);
   adder_mem_array_reg_1_15_inst : dff_asyncrsthl port map( d => N54, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_15_port);
   adder_mem_array_reg_1_16_inst : dff_asyncrsthl port map( d => N55, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_16_port);
   adder_mem_array_reg_1_17_inst : dff_asyncrsthl port map( d => N56, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_17_port);
   adder_mem_array_reg_1_18_inst : dff_asyncrsthl port map( d => N57, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_18_port);
   adder_mem_array_reg_1_19_inst : dff_asyncrsthl port map( d => N58, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_19_port);
   adder_mem_array_reg_1_20_inst : dff_asyncrsthl port map( d => N59, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_20_port);
   adder_mem_array_reg_1_21_inst : dff_asyncrsthl port map( d => N60, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_21_port);
   adder_mem_array_reg_1_22_inst : dff_asyncrsthl port map( d => N61, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_22_port);
   adder_mem_array_reg_1_23_inst : dff_asyncrsthl port map( d => N62, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_23_port);
   adder_mem_array_reg_1_24_inst : dff_asyncrsthl port map( d => N63, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_24_port);
   adder_mem_array_reg_1_25_inst : dff_asyncrsthl port map( d => N64, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_25_port);
   adder_mem_array_reg_1_26_inst : dff_asyncrsthl port map( d => N65, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_26_port);
   adder_mem_array_reg_1_27_inst : dff_asyncrsthl port map( d => N66, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_27_port);
   adder_mem_array_reg_1_28_inst : dff_asyncrsthl port map( d => N67, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_28_port);
   adder_mem_array_reg_1_29_inst : dff_asyncrsthl port map( d => N68, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_29_port);
   adder_mem_array_reg_1_30_inst : dff_asyncrsthl port map( d => N69, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_30_port);
   adder_mem_array_reg_1_31_inst : dff_asyncrsthl port map( d => N70, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_31_port);
   adder_mem_array_reg_1_32_inst : dff_asyncrsthl port map( d => N71, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_1_32_port);
   adder_mem_array_reg_0_0_inst : dff_asyncrsthl port map( d => N6, gclk => clk
                           , asyncrsthl => rst, q => adder_mem_array_0_0_port);
   adder_mem_array_reg_0_1_inst : dff_asyncrsthl port map( d => N7, gclk => clk
                           , asyncrsthl => rst, q => adder_mem_array_0_1_port);
   adder_mem_array_reg_0_2_inst : dff_asyncrsthl port map( d => N8, gclk => clk
                           , asyncrsthl => rst, q => adder_mem_array_0_2_port);
   adder_mem_array_reg_0_3_inst : dff_asyncrsthl port map( d => N9, gclk => clk
                           , asyncrsthl => rst, q => adder_mem_array_0_3_port);
   adder_mem_array_reg_0_4_inst : dff_asyncrsthl port map( d => N10, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_4_port);
   adder_mem_array_reg_0_5_inst : dff_asyncrsthl port map( d => N11, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_5_port);
   adder_mem_array_reg_0_6_inst : dff_asyncrsthl port map( d => N12, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_6_port);
   adder_mem_array_reg_0_7_inst : dff_asyncrsthl port map( d => N13, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_7_port);
   adder_mem_array_reg_0_8_inst : dff_asyncrsthl port map( d => N14, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_8_port);
   adder_mem_array_reg_0_9_inst : dff_asyncrsthl port map( d => N15, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_9_port);
   adder_mem_array_reg_0_10_inst : dff_asyncrsthl port map( d => N16, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_10_port);
   adder_mem_array_reg_0_11_inst : dff_asyncrsthl port map( d => N17, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_11_port);
   adder_mem_array_reg_0_12_inst : dff_asyncrsthl port map( d => N18, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_12_port);
   adder_mem_array_reg_0_13_inst : dff_asyncrsthl port map( d => N19, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_13_port);
   adder_mem_array_reg_0_14_inst : dff_asyncrsthl port map( d => N20, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_14_port);
   adder_mem_array_reg_0_15_inst : dff_asyncrsthl port map( d => N21, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_15_port);
   adder_mem_array_reg_0_16_inst : dff_asyncrsthl port map( d => N22, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_16_port);
   adder_mem_array_reg_0_17_inst : dff_asyncrsthl port map( d => N23, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_17_port);
   adder_mem_array_reg_0_18_inst : dff_asyncrsthl port map( d => N24, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_18_port);
   adder_mem_array_reg_0_19_inst : dff_asyncrsthl port map( d => N25, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_19_port);
   adder_mem_array_reg_0_20_inst : dff_asyncrsthl port map( d => N26, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_20_port);
   adder_mem_array_reg_0_21_inst : dff_asyncrsthl port map( d => N27, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_21_port);
   adder_mem_array_reg_0_22_inst : dff_asyncrsthl port map( d => N28, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_22_port);
   adder_mem_array_reg_0_23_inst : dff_asyncrsthl port map( d => N29, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_23_port);
   adder_mem_array_reg_0_24_inst : dff_asyncrsthl port map( d => N30, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_24_port);
   adder_mem_array_reg_0_25_inst : dff_asyncrsthl port map( d => N31, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_25_port);
   adder_mem_array_reg_0_26_inst : dff_asyncrsthl port map( d => N32, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_26_port);
   adder_mem_array_reg_0_27_inst : dff_asyncrsthl port map( d => N33, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_27_port);
   adder_mem_array_reg_0_28_inst : dff_asyncrsthl port map( d => N34, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_28_port);
   adder_mem_array_reg_0_29_inst : dff_asyncrsthl port map( d => N35, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_29_port);
   adder_mem_array_reg_0_30_inst : dff_asyncrsthl port map( d => N36, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_30_port);
   adder_mem_array_reg_0_31_inst : dff_asyncrsthl port map( d => N37, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_31_port);
   adder_mem_array_reg_0_32_inst : dff_asyncrsthl port map( d => N38, gclk => 
                           clk, asyncrsthl => rst, q => 
                           adder_mem_array_0_32_port);
   coeff_cnt_reg_0_inst : dff port map( d => n206, gclk => clk, rnot => n121, q
                           => coeff_cnt_0_port);
   ready_h_out_reg_reg : dff_asyncprehh port map( d => n205, gclk => clk, 
                           asyncprehh => rst, q => ready_h_out_port);
   coeff_cnt_reg_1_inst : dff port map( d => n204, gclk => clk, rnot => n121, q
                           => coeff_cnt_1_port);
   coefficient_mem_array_reg_3_0_inst : dff port map( d => n203, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_0_port);
   coefficient_mem_array_reg_2_0_inst : dff port map( d => n202, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_0_port);
   coefficient_mem_array_reg_1_0_inst : dff port map( d => n201, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_0_port);
   coefficient_mem_array_reg_0_0_inst : dff port map( d => n200, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_0_port);
   coefficient_mem_array_reg_3_15_inst : dff port map( d => n199, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_15_port);
   coefficient_mem_array_reg_2_15_inst : dff port map( d => n198, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_15_port);
   coefficient_mem_array_reg_1_15_inst : dff port map( d => n197, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_15_port);
   coefficient_mem_array_reg_0_15_inst : dff port map( d => n196, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_15_port);
   coefficient_mem_array_reg_3_14_inst : dff port map( d => n195, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_14_port);
   coefficient_mem_array_reg_2_14_inst : dff port map( d => n194, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_14_port);
   coefficient_mem_array_reg_1_14_inst : dff port map( d => n193, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_14_port);
   coefficient_mem_array_reg_0_14_inst : dff port map( d => n192, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_14_port);
   coefficient_mem_array_reg_3_13_inst : dff port map( d => n191, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_13_port);
   coefficient_mem_array_reg_2_13_inst : dff port map( d => n190, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_13_port);
   coefficient_mem_array_reg_1_13_inst : dff port map( d => n189, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_13_port);
   coefficient_mem_array_reg_0_13_inst : dff port map( d => n188, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_13_port);
   coefficient_mem_array_reg_3_12_inst : dff port map( d => n187, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_12_port);
   coefficient_mem_array_reg_2_12_inst : dff port map( d => n186, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_12_port);
   coefficient_mem_array_reg_1_12_inst : dff port map( d => n185, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_12_port);
   coefficient_mem_array_reg_0_12_inst : dff port map( d => n184, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_12_port);
   coefficient_mem_array_reg_3_11_inst : dff port map( d => n183, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_11_port);
   coefficient_mem_array_reg_2_11_inst : dff port map( d => n182, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_11_port);
   coefficient_mem_array_reg_1_11_inst : dff port map( d => n181, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_11_port);
   coefficient_mem_array_reg_0_11_inst : dff port map( d => n180, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_11_port);
   coefficient_mem_array_reg_3_10_inst : dff port map( d => n179, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_10_port);
   coefficient_mem_array_reg_2_10_inst : dff port map( d => n178, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_10_port);
   coefficient_mem_array_reg_1_10_inst : dff port map( d => n177, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_10_port);
   coefficient_mem_array_reg_0_10_inst : dff port map( d => n176, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_10_port);
   coefficient_mem_array_reg_3_9_inst : dff port map( d => n175, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_9_port);
   coefficient_mem_array_reg_2_9_inst : dff port map( d => n174, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_9_port);
   coefficient_mem_array_reg_1_9_inst : dff port map( d => n173, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_9_port);
   coefficient_mem_array_reg_0_9_inst : dff port map( d => n172, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_9_port);
   coefficient_mem_array_reg_3_8_inst : dff port map( d => n171, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_8_port);
   coefficient_mem_array_reg_2_8_inst : dff port map( d => n170, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_8_port);
   coefficient_mem_array_reg_1_8_inst : dff port map( d => n169, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_8_port);
   coefficient_mem_array_reg_0_8_inst : dff port map( d => n168, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_8_port);
   coefficient_mem_array_reg_3_7_inst : dff port map( d => n167, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_7_port);
   coefficient_mem_array_reg_2_7_inst : dff port map( d => n166, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_7_port);
   coefficient_mem_array_reg_1_7_inst : dff port map( d => n165, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_7_port);
   coefficient_mem_array_reg_0_7_inst : dff port map( d => n164, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_7_port);
   coefficient_mem_array_reg_3_6_inst : dff port map( d => n163, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_6_port);
   coefficient_mem_array_reg_2_6_inst : dff port map( d => n162, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_6_port);
   coefficient_mem_array_reg_1_6_inst : dff port map( d => n161, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_6_port);
   coefficient_mem_array_reg_0_6_inst : dff port map( d => n160, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_6_port);
   coefficient_mem_array_reg_3_5_inst : dff port map( d => n159, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_5_port);
   coefficient_mem_array_reg_2_5_inst : dff port map( d => n158, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_5_port);
   coefficient_mem_array_reg_1_5_inst : dff port map( d => n157, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_5_port);
   coefficient_mem_array_reg_0_5_inst : dff port map( d => n156, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_5_port);
   coefficient_mem_array_reg_3_4_inst : dff port map( d => n155, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_4_port);
   coefficient_mem_array_reg_2_4_inst : dff port map( d => n154, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_4_port);
   coefficient_mem_array_reg_1_4_inst : dff port map( d => n153, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_4_port);
   coefficient_mem_array_reg_0_4_inst : dff port map( d => n152, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_4_port);
   coefficient_mem_array_reg_3_3_inst : dff port map( d => n151, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_3_port);
   coefficient_mem_array_reg_2_3_inst : dff port map( d => n150, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_3_port);
   coefficient_mem_array_reg_1_3_inst : dff port map( d => n149, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_3_port);
   coefficient_mem_array_reg_0_3_inst : dff port map( d => n148, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_3_port);
   coefficient_mem_array_reg_3_2_inst : dff port map( d => n147, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_2_port);
   coefficient_mem_array_reg_2_2_inst : dff port map( d => n146, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_2_port);
   coefficient_mem_array_reg_1_2_inst : dff port map( d => n145, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_2_port);
   coefficient_mem_array_reg_0_2_inst : dff port map( d => n144, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_2_port);
   coefficient_mem_array_reg_3_1_inst : dff port map( d => n143, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_3_1_port);
   coefficient_mem_array_reg_2_1_inst : dff port map( d => n142, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_2_1_port);
   coefficient_mem_array_reg_1_1_inst : dff port map( d => n141, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_1_1_port);
   coefficient_mem_array_reg_0_1_inst : dff port map( d => n140, gclk => clk, 
                           rnot => n121, q => coefficient_mem_array_0_1_port);
   valid_out_reg_reg : dff port map( d => n139, gclk => clk, rnot => n121, q =>
                           valid_out_port);
   ready_x_out_reg_reg : dff port map( d => n138, gclk => clk, rnot => n121, q 
                           => ready_x_out_port);
   input_sample_mem_reg_0_inst : dff port map( d => n137, gclk => clk, rnot => 
                           n121, q => input_sample_mem_0_port);
   input_sample_mem_reg_15_inst : dff port map( d => n136, gclk => clk, rnot =>
                           n121, q => input_sample_mem_15_port);
   input_sample_mem_reg_14_inst : dff port map( d => n135, gclk => clk, rnot =>
                           n121, q => input_sample_mem_14_port);
   input_sample_mem_reg_13_inst : dff port map( d => n134, gclk => clk, rnot =>
                           n121, q => input_sample_mem_13_port);
   input_sample_mem_reg_12_inst : dff port map( d => n133, gclk => clk, rnot =>
                           n121, q => input_sample_mem_12_port);
   input_sample_mem_reg_11_inst : dff port map( d => n132, gclk => clk, rnot =>
                           n121, q => input_sample_mem_11_port);
   input_sample_mem_reg_10_inst : dff port map( d => n131, gclk => clk, rnot =>
                           n121, q => input_sample_mem_10_port);
   input_sample_mem_reg_9_inst : dff port map( d => n130, gclk => clk, rnot => 
                           n121, q => input_sample_mem_9_port);
   input_sample_mem_reg_8_inst : dff port map( d => n129, gclk => clk, rnot => 
                           n121, q => input_sample_mem_8_port);
   input_sample_mem_reg_7_inst : dff port map( d => n128, gclk => clk, rnot => 
                           n121, q => input_sample_mem_7_port);
   input_sample_mem_reg_6_inst : dff port map( d => n127, gclk => clk, rnot => 
                           n121, q => input_sample_mem_6_port);
   input_sample_mem_reg_5_inst : dff port map( d => n126, gclk => clk, rnot => 
                           n121, q => input_sample_mem_5_port);
   input_sample_mem_reg_4_inst : dff port map( d => n125, gclk => clk, rnot => 
                           n121, q => input_sample_mem_4_port);
   input_sample_mem_reg_3_inst : dff port map( d => n124, gclk => clk, rnot => 
                           n121, q => input_sample_mem_3_port);
   input_sample_mem_reg_2_inst : dff port map( d => n123, gclk => clk, rnot => 
                           n121, q => input_sample_mem_2_port);
   input_sample_mem_reg_1_inst : dff port map( d => n122, gclk => clk, rnot => 
                           n121, q => input_sample_mem_1_port);
   U3 : inv port map( inb => n16_port, outb => n139);
   U4 : aoi12 port map( b => coeff_cnt_0_port, c => coeff_cnt_1_port, a => 
                           valid_out_port, outb => n16_port);
   U12 : inv port map( inb => n17_port, outb => n138);
   U13 : aoi12 port map( b => coeff_cnt_0_port, c => coeff_cnt_1_port, a => 
                           ready_x_out_port, outb => n17_port);
   U14 : aoi12 port map( b => coeff_cnt_1_port, c => coeff_cnt_0_port, a => 
                           n18_port, outb => n205);
   U15 : inv port map( inb => ready_h_out_port, outb => n18_port);
   U16 : inv port map( inb => n19_port, outb => n130);
   U17 : aoi22 port map( a => x_data_in(9), b => n20_port, c => 
                           input_sample_mem_9_port, d => n21_port, outb => 
                           n19_port);
   U18 : inv port map( inb => n22_port, outb => n129);
   U19 : aoi22 port map( a => x_data_in(8), b => n20_port, c => 
                           input_sample_mem_8_port, d => n21_port, outb => 
                           n22_port);
   U20 : inv port map( inb => n23_port, outb => n128);
   U21 : aoi22 port map( a => x_data_in(7), b => n20_port, c => 
                           input_sample_mem_7_port, d => n21_port, outb => 
                           n23_port);
   U22 : inv port map( inb => n24_port, outb => n127);
   U23 : aoi22 port map( a => x_data_in(6), b => n20_port, c => 
                           input_sample_mem_6_port, d => n21_port, outb => 
                           n24_port);
   U24 : inv port map( inb => n25_port, outb => n126);
   U25 : aoi22 port map( a => x_data_in(5), b => n20_port, c => 
                           input_sample_mem_5_port, d => n21_port, outb => 
                           n25_port);
   U26 : inv port map( inb => n26_port, outb => n125);
   U27 : aoi22 port map( a => x_data_in(4), b => n20_port, c => 
                           input_sample_mem_4_port, d => n21_port, outb => 
                           n26_port);
   U28 : inv port map( inb => n27_port, outb => n124);
   U29 : aoi22 port map( a => x_data_in(3), b => n20_port, c => 
                           input_sample_mem_3_port, d => n21_port, outb => 
                           n27_port);
   U30 : inv port map( inb => n28_port, outb => n123);
   U31 : aoi22 port map( a => x_data_in(2), b => n20_port, c => 
                           input_sample_mem_2_port, d => n21_port, outb => 
                           n28_port);
   U32 : inv port map( inb => n29_port, outb => n122);
   U33 : aoi22 port map( a => x_data_in(1), b => n20_port, c => 
                           input_sample_mem_1_port, d => n21_port, outb => 
                           n29_port);
   U34 : inv port map( inb => n30_port, outb => n136);
   U35 : aoi22 port map( a => x_data_in(15), b => n20_port, c => 
                           input_sample_mem_15_port, d => n21_port, outb => 
                           n30_port);
   U36 : inv port map( inb => n31_port, outb => n135);
   U37 : aoi22 port map( a => x_data_in(14), b => n20_port, c => 
                           input_sample_mem_14_port, d => n21_port, outb => 
                           n31_port);
   U38 : inv port map( inb => n32_port, outb => n134);
   U39 : aoi22 port map( a => x_data_in(13), b => n20_port, c => 
                           input_sample_mem_13_port, d => n21_port, outb => 
                           n32_port);
   U40 : inv port map( inb => n33_port, outb => n133);
   U41 : aoi22 port map( a => x_data_in(12), b => n20_port, c => 
                           input_sample_mem_12_port, d => n21_port, outb => 
                           n33_port);
   U42 : inv port map( inb => n34_port, outb => n132);
   U43 : aoi22 port map( a => x_data_in(11), b => n20_port, c => 
                           input_sample_mem_11_port, d => n21_port, outb => 
                           n34_port);
   U44 : inv port map( inb => n35_port, outb => n131);
   U45 : aoi22 port map( a => x_data_in(10), b => n20_port, c => 
                           input_sample_mem_10_port, d => n21_port, outb => 
                           n35_port);
   U46 : inv port map( inb => n36_port, outb => n137);
   U47 : aoi22 port map( a => x_data_in(0), b => n20_port, c => 
                           input_sample_mem_0_port, d => n21_port, outb => 
                           n36_port);
   U48 : inv port map( inb => n21_port, outb => n20_port);
   U49 : nand2 port map( a => valid_x_in, b => ready_x_out_port, outb => 
                           n21_port);
   U50 : inv port map( inb => n37_port, outb => n175);
   U51 : aoi22 port map( a => n38_port, b => h_data_in(9), c => n39_port, d => 
                           coefficient_mem_array_3_9_port, outb => n37_port);
   U52 : inv port map( inb => n40_port, outb => n171);
   U53 : aoi22 port map( a => n38_port, b => h_data_in(8), c => n39_port, d => 
                           coefficient_mem_array_3_8_port, outb => n40_port);
   U54 : inv port map( inb => n41_port, outb => n167);
   U55 : aoi22 port map( a => n38_port, b => h_data_in(7), c => n39_port, d => 
                           coefficient_mem_array_3_7_port, outb => n41_port);
   U56 : inv port map( inb => n42_port, outb => n163);
   U57 : aoi22 port map( a => n38_port, b => h_data_in(6), c => n39_port, d => 
                           coefficient_mem_array_3_6_port, outb => n42_port);
   U58 : inv port map( inb => n43_port, outb => n159);
   U59 : aoi22 port map( a => n38_port, b => h_data_in(5), c => n39_port, d => 
                           coefficient_mem_array_3_5_port, outb => n43_port);
   U60 : inv port map( inb => n44_port, outb => n155);
   U61 : aoi22 port map( a => n38_port, b => h_data_in(4), c => n39_port, d => 
                           coefficient_mem_array_3_4_port, outb => n44_port);
   U62 : inv port map( inb => n45_port, outb => n151);
   U63 : aoi22 port map( a => n38_port, b => h_data_in(3), c => n39_port, d => 
                           coefficient_mem_array_3_3_port, outb => n45_port);
   U64 : inv port map( inb => n46_port, outb => n147);
   U65 : aoi22 port map( a => n38_port, b => h_data_in(2), c => n39_port, d => 
                           coefficient_mem_array_3_2_port, outb => n46_port);
   U66 : inv port map( inb => n47_port, outb => n143);
   U67 : aoi22 port map( a => n38_port, b => h_data_in(1), c => n39_port, d => 
                           coefficient_mem_array_3_1_port, outb => n47_port);
   U68 : inv port map( inb => n48_port, outb => n199);
   U69 : aoi22 port map( a => n38_port, b => h_data_in(15), c => n39_port, d =>
                           coefficient_mem_array_3_15_port, outb => n48_port);
   U70 : inv port map( inb => n49_port, outb => n195);
   U71 : aoi22 port map( a => n38_port, b => h_data_in(14), c => n39_port, d =>
                           coefficient_mem_array_3_14_port, outb => n49_port);
   U72 : inv port map( inb => n50_port, outb => n191);
   U73 : aoi22 port map( a => n38_port, b => h_data_in(13), c => n39_port, d =>
                           coefficient_mem_array_3_13_port, outb => n50_port);
   U74 : inv port map( inb => n51_port, outb => n187);
   U75 : aoi22 port map( a => n38_port, b => h_data_in(12), c => n39_port, d =>
                           coefficient_mem_array_3_12_port, outb => n51_port);
   U76 : inv port map( inb => n52_port, outb => n183);
   U77 : aoi22 port map( a => n38_port, b => h_data_in(11), c => n39_port, d =>
                           coefficient_mem_array_3_11_port, outb => n52_port);
   U78 : inv port map( inb => n53_port, outb => n179);
   U79 : aoi22 port map( a => n38_port, b => h_data_in(10), c => n39_port, d =>
                           coefficient_mem_array_3_10_port, outb => n53_port);
   U80 : inv port map( inb => n54_port, outb => n203);
   U81 : aoi22 port map( a => n38_port, b => h_data_in(0), c => n39_port, d => 
                           coefficient_mem_array_3_0_port, outb => n54_port);
   U82 : oai22 port map( a => n55_port, b => n39_port, c => n38_port, d => 
                           n56_port, outb => n174);
   U83 : inv port map( inb => coefficient_mem_array_3_9_port, outb => n55_port)
                           ;
   U84 : oai22 port map( a => n39_port, b => n57_port, c => n38_port, d => 
                           n58_port, outb => n170);
   U85 : inv port map( inb => coefficient_mem_array_3_8_port, outb => n57_port)
                           ;
   U86 : oai22 port map( a => n39_port, b => n59_port, c => n38_port, d => 
                           n60_port, outb => n166);
   U87 : inv port map( inb => coefficient_mem_array_3_7_port, outb => n59_port)
                           ;
   U88 : oai22 port map( a => n39_port, b => n61_port, c => n38_port, d => 
                           n62_port, outb => n162);
   U89 : inv port map( inb => coefficient_mem_array_3_6_port, outb => n61_port)
                           ;
   U90 : oai22 port map( a => n39_port, b => n63_port, c => n38_port, d => 
                           n64_port, outb => n158);
   U91 : inv port map( inb => coefficient_mem_array_3_5_port, outb => n63_port)
                           ;
   U92 : oai22 port map( a => n39_port, b => n65_port, c => n38_port, d => 
                           n66_port, outb => n154);
   U93 : inv port map( inb => coefficient_mem_array_3_4_port, outb => n65_port)
                           ;
   U94 : oai22 port map( a => n39_port, b => n67_port, c => n38_port, d => 
                           n68_port, outb => n150);
   U95 : inv port map( inb => coefficient_mem_array_3_3_port, outb => n67_port)
                           ;
   U96 : oai22 port map( a => n39_port, b => n69_port, c => n38_port, d => 
                           n70_port, outb => n146);
   U97 : inv port map( inb => coefficient_mem_array_3_2_port, outb => n69_port)
                           ;
   U98 : oai22 port map( a => n39_port, b => n71_port, c => n38_port, d => 
                           n72_port, outb => n142);
   U99 : inv port map( inb => coefficient_mem_array_3_1_port, outb => n71_port)
                           ;
   U100 : oai22 port map( a => n39_port, b => n73_port, c => n38_port, d => 
                           n74_port, outb => n198);
   U101 : inv port map( inb => coefficient_mem_array_3_15_port, outb => 
                           n73_port);
   U102 : oai22 port map( a => n39_port, b => n75_port, c => n38_port, d => 
                           n76_port, outb => n194);
   U103 : inv port map( inb => coefficient_mem_array_3_14_port, outb => 
                           n75_port);
   U104 : oai22 port map( a => n39_port, b => n77_port, c => n38_port, d => 
                           n78_port, outb => n190);
   U105 : inv port map( inb => coefficient_mem_array_3_13_port, outb => 
                           n77_port);
   U106 : oai22 port map( a => n39_port, b => n79_port, c => n38_port, d => 
                           n80_port, outb => n186);
   U107 : inv port map( inb => coefficient_mem_array_3_12_port, outb => 
                           n79_port);
   U108 : oai22 port map( a => n39_port, b => n81_port, c => n38_port, d => 
                           n82_port, outb => n182);
   U109 : inv port map( inb => coefficient_mem_array_3_11_port, outb => 
                           n81_port);
   U110 : oai22 port map( a => n39_port, b => n83_port, c => n38_port, d => 
                           n84_port, outb => n178);
   U111 : inv port map( inb => coefficient_mem_array_3_10_port, outb => 
                           n83_port);
   U112 : oai22 port map( a => n39_port, b => n85_port, c => n38_port, d => 
                           n86_port, outb => n202);
   U113 : inv port map( inb => coefficient_mem_array_3_0_port, outb => n85_port
                           );
   U114 : oai22 port map( a => n39_port, b => n56_port, c => n38_port, d => 
                           n87_port, outb => n173);
   U115 : inv port map( inb => coefficient_mem_array_2_9_port, outb => n56_port
                           );
   U116 : oai22 port map( a => n39_port, b => n58_port, c => n38_port, d => 
                           n88_port, outb => n169);
   U117 : inv port map( inb => coefficient_mem_array_2_8_port, outb => n58_port
                           );
   U118 : oai22 port map( a => n39_port, b => n60_port, c => n38_port, d => 
                           n89_port, outb => n165);
   U119 : inv port map( inb => coefficient_mem_array_2_7_port, outb => n60_port
                           );
   U120 : oai22 port map( a => n39_port, b => n62_port, c => n38_port, d => 
                           n90_port, outb => n161);
   U121 : inv port map( inb => coefficient_mem_array_2_6_port, outb => n62_port
                           );
   U122 : oai22 port map( a => n39_port, b => n64_port, c => n38_port, d => 
                           n91_port, outb => n157);
   U123 : inv port map( inb => coefficient_mem_array_2_5_port, outb => n64_port
                           );
   U124 : oai22 port map( a => n39_port, b => n66_port, c => n38_port, d => 
                           n92_port, outb => n153);
   U125 : inv port map( inb => coefficient_mem_array_2_4_port, outb => n66_port
                           );
   U126 : oai22 port map( a => n39_port, b => n68_port, c => n38_port, d => 
                           n93_port, outb => n149);
   U127 : inv port map( inb => coefficient_mem_array_2_3_port, outb => n68_port
                           );
   U128 : oai22 port map( a => n39_port, b => n70_port, c => n38_port, d => 
                           n94_port, outb => n145);
   U129 : inv port map( inb => coefficient_mem_array_2_2_port, outb => n70_port
                           );
   U130 : oai22 port map( a => n39_port, b => n72_port, c => n38_port, d => 
                           n95_port, outb => n141);
   U131 : inv port map( inb => coefficient_mem_array_2_1_port, outb => n72_port
                           );
   U132 : oai22 port map( a => n39_port, b => n74_port, c => n38_port, d => 
                           n96_port, outb => n197);
   U133 : inv port map( inb => coefficient_mem_array_2_15_port, outb => 
                           n74_port);
   U134 : oai22 port map( a => n39_port, b => n76_port, c => n38_port, d => 
                           n97_port, outb => n193);
   U135 : inv port map( inb => coefficient_mem_array_2_14_port, outb => 
                           n76_port);
   U136 : oai22 port map( a => n39_port, b => n78_port, c => n38_port, d => 
                           n98_port, outb => n189);
   U137 : inv port map( inb => coefficient_mem_array_2_13_port, outb => 
                           n78_port);
   U138 : oai22 port map( a => n39_port, b => n80_port, c => n38_port, d => 
                           n99_port, outb => n185);
   U139 : inv port map( inb => coefficient_mem_array_2_12_port, outb => 
                           n80_port);
   U140 : oai22 port map( a => n39_port, b => n82_port, c => n38_port, d => 
                           n100_port, outb => n181);
   U141 : inv port map( inb => coefficient_mem_array_2_11_port, outb => 
                           n82_port);
   U142 : oai22 port map( a => n39_port, b => n84_port, c => n38_port, d => 
                           n101_port, outb => n177);
   U143 : inv port map( inb => coefficient_mem_array_2_10_port, outb => 
                           n84_port);
   U144 : oai22 port map( a => n39_port, b => n86_port, c => n38_port, d => 
                           n102_port, outb => n201);
   U145 : inv port map( inb => coefficient_mem_array_2_0_port, outb => n86_port
                           );
   U146 : oai12 port map( b => n39_port, c => n87_port, a => n103_port, outb =>
                           n172);
   U147 : nand2 port map( a => coefficient_mem_array_0_9_port, b => n39_port, 
                           outb => n103_port);
   U148 : inv port map( inb => coefficient_mem_array_1_9_port, outb => n87_port
                           );
   U149 : oai12 port map( b => n39_port, c => n88_port, a => n104_port, outb =>
                           n168);
   U150 : nand2 port map( a => coefficient_mem_array_0_8_port, b => n39_port, 
                           outb => n104_port);
   U151 : inv port map( inb => coefficient_mem_array_1_8_port, outb => n88_port
                           );
   U152 : oai12 port map( b => n39_port, c => n89_port, a => n105, outb => n164
                           );
   U153 : nand2 port map( a => coefficient_mem_array_0_7_port, b => n39_port, 
                           outb => n105);
   U154 : inv port map( inb => coefficient_mem_array_1_7_port, outb => n89_port
                           );
   U155 : oai12 port map( b => n39_port, c => n90_port, a => n106, outb => n160
                           );
   U156 : nand2 port map( a => coefficient_mem_array_0_6_port, b => n39_port, 
                           outb => n106);
   U157 : inv port map( inb => coefficient_mem_array_1_6_port, outb => n90_port
                           );
   U158 : oai12 port map( b => n39_port, c => n91_port, a => n107, outb => n156
                           );
   U159 : nand2 port map( a => coefficient_mem_array_0_5_port, b => n39_port, 
                           outb => n107);
   U160 : inv port map( inb => coefficient_mem_array_1_5_port, outb => n91_port
                           );
   U161 : oai12 port map( b => n39_port, c => n92_port, a => n108, outb => n152
                           );
   U162 : nand2 port map( a => coefficient_mem_array_0_4_port, b => n39_port, 
                           outb => n108);
   U163 : inv port map( inb => coefficient_mem_array_1_4_port, outb => n92_port
                           );
   U164 : oai12 port map( b => n39_port, c => n93_port, a => n109, outb => n148
                           );
   U165 : nand2 port map( a => coefficient_mem_array_0_3_port, b => n39_port, 
                           outb => n109);
   U166 : inv port map( inb => coefficient_mem_array_1_3_port, outb => n93_port
                           );
   U167 : oai12 port map( b => n39_port, c => n94_port, a => n110, outb => n144
                           );
   U168 : nand2 port map( a => coefficient_mem_array_0_2_port, b => n39_port, 
                           outb => n110);
   U169 : inv port map( inb => coefficient_mem_array_1_2_port, outb => n94_port
                           );
   U170 : oai12 port map( b => n39_port, c => n95_port, a => n111, outb => n140
                           );
   U171 : nand2 port map( a => coefficient_mem_array_0_1_port, b => n39_port, 
                           outb => n111);
   U172 : inv port map( inb => coefficient_mem_array_1_1_port, outb => n95_port
                           );
   U173 : oai12 port map( b => n39_port, c => n96_port, a => n112, outb => n196
                           );
   U174 : nand2 port map( a => coefficient_mem_array_0_15_port, b => n39_port, 
                           outb => n112);
   U175 : inv port map( inb => coefficient_mem_array_1_15_port, outb => 
                           n96_port);
   U176 : oai12 port map( b => n39_port, c => n97_port, a => n113, outb => n192
                           );
   U177 : nand2 port map( a => coefficient_mem_array_0_14_port, b => n39_port, 
                           outb => n113);
   U178 : inv port map( inb => coefficient_mem_array_1_14_port, outb => 
                           n97_port);
   U179 : oai12 port map( b => n39_port, c => n98_port, a => n114, outb => n188
                           );
   U180 : nand2 port map( a => coefficient_mem_array_0_13_port, b => n39_port, 
                           outb => n114);
   U181 : inv port map( inb => coefficient_mem_array_1_13_port, outb => 
                           n98_port);
   U182 : oai12 port map( b => n39_port, c => n99_port, a => n115, outb => n184
                           );
   U183 : nand2 port map( a => coefficient_mem_array_0_12_port, b => n39_port, 
                           outb => n115);
   U184 : inv port map( inb => coefficient_mem_array_1_12_port, outb => 
                           n99_port);
   U185 : oai12 port map( b => n39_port, c => n100_port, a => n116, outb => 
                           n180);
   U186 : nand2 port map( a => coefficient_mem_array_0_11_port, b => n39_port, 
                           outb => n116);
   U187 : inv port map( inb => coefficient_mem_array_1_11_port, outb => 
                           n100_port);
   U188 : oai12 port map( b => n39_port, c => n101_port, a => n117, outb => 
                           n176);
   U189 : nand2 port map( a => coefficient_mem_array_0_10_port, b => n39_port, 
                           outb => n117);
   U190 : inv port map( inb => coefficient_mem_array_1_10_port, outb => 
                           n101_port);
   U191 : oai12 port map( b => n39_port, c => n102_port, a => n118, outb => 
                           n200);
   U192 : nand2 port map( a => coefficient_mem_array_0_0_port, b => n39_port, 
                           outb => n118);
   U193 : inv port map( inb => coefficient_mem_array_1_0_port, outb => 
                           n102_port);
   U194 : xor2 port map( a => n119, b => n120, outb => n204);
   U195 : nand2 port map( a => coeff_cnt_0_port, b => n38_port, outb => n120);
   U196 : inv port map( inb => coeff_cnt_1_port, outb => n119);
   U197 : inv port map( inb => rst, outb => n121);
   U198 : xor2 port map( a => coeff_cnt_0_port, b => n38_port, outb => n206);
   U199 : inv port map( inb => n39_port, outb => n38_port);
   U200 : nand2 port map( a => valid_h_in, b => ready_h_out_port, outb => 
                           n39_port);
   U201 : inv port map( inb => n207, outb => y_data_out(9));
   U202 : nand2 port map( a => valid_out_port, b => adder_mem_array_0_9_port, 
                           outb => n207);
   U203 : inv port map( inb => n208, outb => y_data_out(8));
   U204 : nand2 port map( a => adder_mem_array_0_8_port, b => valid_out_port, 
                           outb => n208);
   U205 : inv port map( inb => n209, outb => y_data_out(7));
   U206 : nand2 port map( a => adder_mem_array_0_7_port, b => valid_out_port, 
                           outb => n209);
   U207 : inv port map( inb => n210, outb => y_data_out(6));
   U208 : nand2 port map( a => adder_mem_array_0_6_port, b => valid_out_port, 
                           outb => n210);
   U209 : inv port map( inb => n211, outb => y_data_out(5));
   U210 : nand2 port map( a => adder_mem_array_0_5_port, b => valid_out_port, 
                           outb => n211);
   U211 : inv port map( inb => n212, outb => y_data_out(4));
   U212 : nand2 port map( a => adder_mem_array_0_4_port, b => valid_out_port, 
                           outb => n212);
   U213 : inv port map( inb => n213, outb => y_data_out(3));
   U214 : nand2 port map( a => adder_mem_array_0_3_port, b => valid_out_port, 
                           outb => n213);
   U215 : inv port map( inb => n214, outb => y_data_out(32));
   U216 : nand2 port map( a => adder_mem_array_0_32_port, b => valid_out_port, 
                           outb => n214);
   U217 : inv port map( inb => n215, outb => y_data_out(31));
   U218 : nand2 port map( a => adder_mem_array_0_31_port, b => valid_out_port, 
                           outb => n215);
   U219 : inv port map( inb => n216, outb => y_data_out(30));
   U220 : nand2 port map( a => adder_mem_array_0_30_port, b => valid_out_port, 
                           outb => n216);
   U221 : inv port map( inb => n217, outb => y_data_out(2));
   U222 : nand2 port map( a => adder_mem_array_0_2_port, b => valid_out_port, 
                           outb => n217);
   U223 : inv port map( inb => n218, outb => y_data_out(29));
   U224 : nand2 port map( a => adder_mem_array_0_29_port, b => valid_out_port, 
                           outb => n218);
   U225 : inv port map( inb => n219, outb => y_data_out(28));
   U226 : nand2 port map( a => adder_mem_array_0_28_port, b => valid_out_port, 
                           outb => n219);
   U227 : inv port map( inb => n220, outb => y_data_out(27));
   U228 : nand2 port map( a => adder_mem_array_0_27_port, b => valid_out_port, 
                           outb => n220);
   U229 : inv port map( inb => n221, outb => y_data_out(26));
   U230 : nand2 port map( a => adder_mem_array_0_26_port, b => valid_out_port, 
                           outb => n221);
   U231 : inv port map( inb => n222, outb => y_data_out(25));
   U232 : nand2 port map( a => adder_mem_array_0_25_port, b => valid_out_port, 
                           outb => n222);
   U233 : inv port map( inb => n223, outb => y_data_out(24));
   U234 : nand2 port map( a => adder_mem_array_0_24_port, b => valid_out_port, 
                           outb => n223);
   U235 : inv port map( inb => n224, outb => y_data_out(23));
   U236 : nand2 port map( a => adder_mem_array_0_23_port, b => valid_out_port, 
                           outb => n224);
   U237 : inv port map( inb => n225, outb => y_data_out(22));
   U238 : nand2 port map( a => adder_mem_array_0_22_port, b => valid_out_port, 
                           outb => n225);
   U239 : inv port map( inb => n226, outb => y_data_out(21));
   U240 : nand2 port map( a => adder_mem_array_0_21_port, b => valid_out_port, 
                           outb => n226);
   U241 : inv port map( inb => n227, outb => y_data_out(20));
   U242 : nand2 port map( a => adder_mem_array_0_20_port, b => valid_out_port, 
                           outb => n227);
   U243 : inv port map( inb => n228, outb => y_data_out(1));
   U244 : nand2 port map( a => adder_mem_array_0_1_port, b => valid_out_port, 
                           outb => n228);
   U245 : inv port map( inb => n229, outb => y_data_out(19));
   U246 : nand2 port map( a => adder_mem_array_0_19_port, b => valid_out_port, 
                           outb => n229);
   U247 : inv port map( inb => n230, outb => y_data_out(18));
   U248 : nand2 port map( a => adder_mem_array_0_18_port, b => valid_out_port, 
                           outb => n230);
   U249 : inv port map( inb => n231, outb => y_data_out(17));
   U250 : nand2 port map( a => adder_mem_array_0_17_port, b => valid_out_port, 
                           outb => n231);
   U251 : inv port map( inb => n232, outb => y_data_out(16));
   U252 : nand2 port map( a => adder_mem_array_0_16_port, b => valid_out_port, 
                           outb => n232);
   U253 : inv port map( inb => n233, outb => y_data_out(15));
   U254 : nand2 port map( a => adder_mem_array_0_15_port, b => valid_out_port, 
                           outb => n233);
   U255 : inv port map( inb => n234, outb => y_data_out(14));
   U256 : nand2 port map( a => adder_mem_array_0_14_port, b => valid_out_port, 
                           outb => n234);
   U257 : inv port map( inb => n235, outb => y_data_out(13));
   U258 : nand2 port map( a => adder_mem_array_0_13_port, b => valid_out_port, 
                           outb => n235);
   U259 : inv port map( inb => n236, outb => y_data_out(12));
   U260 : nand2 port map( a => adder_mem_array_0_12_port, b => valid_out_port, 
                           outb => n236);
   U261 : inv port map( inb => n237, outb => y_data_out(11));
   U262 : nand2 port map( a => adder_mem_array_0_11_port, b => valid_out_port, 
                           outb => n237);
   U263 : inv port map( inb => n238, outb => y_data_out(10));
   U264 : nand2 port map( a => adder_mem_array_0_10_port, b => valid_out_port, 
                           outb => n238);
   U265 : inv port map( inb => n239, outb => y_data_out(0));
   U266 : nand2 port map( a => adder_mem_array_0_0_port, b => valid_out_port, 
                           outb => n239);
   mult_125_G3_FS_1_U6_1_1_3 : oai12 port map( b => n6032, c => n6033, a => 
                           n6034, outb => mult_125_G3_FS_1_C_1_7_0_port);
   mult_125_G3_FS_1_U6_1_1_2 : oai12 port map( b => n6029, c => n6030, a => 
                           n6031, outb => mult_125_G3_FS_1_C_1_6_0_port);
   mult_125_G3_FS_1_U6_1_1_1 : oai12 port map( b => n6026, c => n6027, a => 
                           n6028, outb => mult_125_G3_FS_1_C_1_5_0_port);
   mult_125_G3_FS_1_U6_0_7_1 : oai12 port map( b => n6023, c => n6024, a => 
                           mult_125_G3_FS_1_G_n_int_0_7_0_port, outb => 
                           mult_125_G3_FS_1_C_1_7_1_port);
   mult_125_G3_FS_1_U3_C_0_7_1 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_7_1_port, b => 
                           mult_125_G3_FS_1_C_1_7_1_port, outb => 
                           multiplier_sigs_2_31_port);
   mult_125_G3_FS_1_U3_B_0_7_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_7_1_port, b => 
                           mult_125_G3_FS_1_P_0_7_1_port, outb => n6022);
   mult_125_G3_FS_1_U2_0_7_1 : nand2 port map( a => mult_125_G3_A1_29_port, b 
                           => mult_125_G3_A2_29_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_7_1_port);
   mult_125_G3_FS_1_U1_0_7_1 : nand2 port map( a => n6020, b => n6021, outb => 
                           mult_125_G3_FS_1_P_0_7_1_port);
   mult_125_G3_FS_1_U3_C_0_7_0 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_7_0_port, b => 
                           mult_125_G3_FS_1_C_1_7_0_port, outb => 
                           multiplier_sigs_2_30_port);
   mult_125_G3_FS_1_U3_B_0_7_0 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_7_0_port, b => 
                           mult_125_G3_FS_1_TEMP_P_0_7_0_port, outb => n6019);
   mult_125_G3_FS_1_U2_0_7_0 : nand2 port map( a => mult_125_G3_A1_28_port, b 
                           => mult_125_G3_A2_28_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_7_0_port);
   mult_125_G3_FS_1_U1_0_7_0 : nand2 port map( a => n6017, b => n6018, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_7_0_port);
   mult_125_G3_FS_1_U6_0_6_3 : oai12 port map( b => n6015, c => n6016, a => 
                           mult_125_G3_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G3_FS_1_C_1_6_3_port);
   mult_125_G3_FS_1_U5_0_6_3 : oai12 port map( b => n6013, c => n6014, a => 
                           mult_125_G3_FS_1_G_n_int_0_6_3_port, outb => 
                           mult_125_G3_FS_1_G_1_1_2_port);
   mult_125_G3_FS_1_U4_0_6_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_6_2_port, b => 
                           mult_125_G3_FS_1_P_0_6_3_port, outb => n6033);
   mult_125_G3_FS_1_U3_C_0_6_3 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_6_3_port, b => 
                           mult_125_G3_FS_1_C_1_6_3_port, outb => 
                           multiplier_sigs_2_29_port);
   mult_125_G3_FS_1_U3_B_0_6_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_6_3_port, b => 
                           mult_125_G3_FS_1_P_0_6_3_port, outb => n6012);
   mult_125_G3_FS_1_U2_0_6_3 : nand2 port map( a => mult_125_G3_A1_27_port, b 
                           => mult_125_G3_A2_27_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_6_3_port);
   mult_125_G3_FS_1_U1_0_6_3 : nand2 port map( a => n6010, b => n6011, outb => 
                           mult_125_G3_FS_1_P_0_6_3_port);
   mult_125_G3_FS_1_U6_0_6_2 : oai12 port map( b => n6008, c => n6009, a => 
                           mult_125_G3_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G3_FS_1_C_1_6_2_port);
   mult_125_G3_FS_1_U5_0_6_2 : oai12 port map( b => n6007, c => n6016, a => 
                           mult_125_G3_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_6_2_port);
   mult_125_G3_FS_1_U4_0_6_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_6_1_port, b => 
                           mult_125_G3_FS_1_P_0_6_2_port, outb => n6006);
   mult_125_G3_FS_1_U3_C_0_6_2 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_6_2_port, b => 
                           mult_125_G3_FS_1_C_1_6_2_port, outb => 
                           multiplier_sigs_2_28_port);
   mult_125_G3_FS_1_U3_B_0_6_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_6_2_port, b => 
                           mult_125_G3_FS_1_P_0_6_2_port, outb => n6005);
   mult_125_G3_FS_1_U2_0_6_2 : nand2 port map( a => mult_125_G3_A1_26_port, b 
                           => mult_125_G3_A2_26_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_6_2_port);
   mult_125_G3_FS_1_U1_0_6_2 : nand2 port map( a => n6003, b => n6004, outb => 
                           mult_125_G3_FS_1_P_0_6_2_port);
   mult_125_G3_FS_1_U6_0_6_1 : oai12 port map( b => n6032, c => n6002, a => 
                           mult_125_G3_FS_1_G_n_int_0_6_0_port, outb => 
                           mult_125_G3_FS_1_C_1_6_1_port);
   mult_125_G3_FS_1_U5_0_6_1 : oai12 port map( b => 
                           mult_125_G3_FS_1_G_n_int_0_6_0_port, c => n6009, a 
                           => mult_125_G3_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_6_1_port);
   mult_125_G3_FS_1_U4_0_6_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_6_0_port, b => 
                           mult_125_G3_FS_1_P_0_6_1_port, outb => n6001);
   mult_125_G3_FS_1_U3_C_0_6_1 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_6_1_port, b => 
                           mult_125_G3_FS_1_C_1_6_1_port, outb => 
                           multiplier_sigs_2_27_port);
   mult_125_G3_FS_1_U3_B_0_6_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_6_1_port, b => 
                           mult_125_G3_FS_1_P_0_6_1_port, outb => n6000);
   mult_125_G3_FS_1_U2_0_6_1 : nand2 port map( a => mult_125_G3_A1_25_port, b 
                           => mult_125_G3_A2_25_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_6_1_port);
   mult_125_G3_FS_1_U1_0_6_1 : nand2 port map( a => n5998, b => n5999, outb => 
                           mult_125_G3_FS_1_P_0_6_1_port);
   mult_125_G3_FS_1_U3_C_0_6_0 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_6_0_port, b => 
                           mult_125_G3_FS_1_C_1_6_0_port, outb => 
                           multiplier_sigs_2_26_port);
   mult_125_G3_FS_1_U3_B_0_6_0 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_6_0_port, b => 
                           mult_125_G3_FS_1_TEMP_P_0_6_0_port, outb => n5997);
   mult_125_G3_FS_1_U2_0_6_0 : nand2 port map( a => mult_125_G3_A1_24_port, b 
                           => mult_125_G3_A2_24_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_6_0_port);
   mult_125_G3_FS_1_U1_0_6_0 : nand2 port map( a => n5995, b => n5996, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_6_0_port);
   mult_125_G3_FS_1_U6_0_5_3 : oai12 port map( b => n5993, c => n5994, a => 
                           mult_125_G3_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G3_FS_1_C_1_5_3_port);
   mult_125_G3_FS_1_U5_0_5_3 : oai12 port map( b => n5991, c => n5992, a => 
                           mult_125_G3_FS_1_G_n_int_0_5_3_port, outb => 
                           mult_125_G3_FS_1_G_1_1_1_port);
   mult_125_G3_FS_1_U4_0_5_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_5_2_port, b => 
                           mult_125_G3_FS_1_P_0_5_3_port, outb => n6030);
   mult_125_G3_FS_1_U3_C_0_5_3 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_5_3_port, b => 
                           mult_125_G3_FS_1_C_1_5_3_port, outb => 
                           multiplier_sigs_2_25_port);
   mult_125_G3_FS_1_U3_B_0_5_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_5_3_port, b => 
                           mult_125_G3_FS_1_P_0_5_3_port, outb => n5990);
   mult_125_G3_FS_1_U2_0_5_3 : nand2 port map( a => mult_125_G3_A1_23_port, b 
                           => mult_125_G3_A2_23_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_5_3_port);
   mult_125_G3_FS_1_U1_0_5_3 : nand2 port map( a => n5988, b => n5989, outb => 
                           mult_125_G3_FS_1_P_0_5_3_port);
   mult_125_G3_FS_1_U6_0_5_2 : oai12 port map( b => n5986, c => n5987, a => 
                           mult_125_G3_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G3_FS_1_C_1_5_2_port);
   mult_125_G3_FS_1_U5_0_5_2 : oai12 port map( b => n5985, c => n5994, a => 
                           mult_125_G3_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_5_2_port);
   mult_125_G3_FS_1_U4_0_5_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_5_1_port, b => 
                           mult_125_G3_FS_1_P_0_5_2_port, outb => n5984);
   mult_125_G3_FS_1_U3_C_0_5_2 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_5_2_port, b => 
                           mult_125_G3_FS_1_C_1_5_2_port, outb => 
                           multiplier_sigs_2_24_port);
   mult_125_G3_FS_1_U3_B_0_5_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_5_2_port, b => 
                           mult_125_G3_FS_1_P_0_5_2_port, outb => n5983);
   mult_125_G3_FS_1_U2_0_5_2 : nand2 port map( a => mult_125_G3_A1_22_port, b 
                           => mult_125_G3_A2_22_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_5_2_port);
   mult_125_G3_FS_1_U1_0_5_2 : nand2 port map( a => n5981, b => n5982, outb => 
                           mult_125_G3_FS_1_P_0_5_2_port);
   mult_125_G3_FS_1_U6_0_5_1 : oai12 port map( b => n6029, c => n5980, a => 
                           mult_125_G3_FS_1_G_n_int_0_5_0_port, outb => 
                           mult_125_G3_FS_1_C_1_5_1_port);
   mult_125_G3_FS_1_U5_0_5_1 : oai12 port map( b => 
                           mult_125_G3_FS_1_G_n_int_0_5_0_port, c => n5987, a 
                           => mult_125_G3_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_5_1_port);
   mult_125_G3_FS_1_U4_0_5_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_5_0_port, b => 
                           mult_125_G3_FS_1_P_0_5_1_port, outb => n5979);
   mult_125_G3_FS_1_U3_C_0_5_1 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_5_1_port, b => 
                           mult_125_G3_FS_1_C_1_5_1_port, outb => 
                           multiplier_sigs_2_23_port);
   mult_125_G3_FS_1_U3_B_0_5_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_5_1_port, b => 
                           mult_125_G3_FS_1_P_0_5_1_port, outb => n5978);
   mult_125_G3_FS_1_U2_0_5_1 : nand2 port map( a => mult_125_G3_A1_21_port, b 
                           => mult_125_G3_A2_21_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_5_1_port);
   mult_125_G3_FS_1_U1_0_5_1 : nand2 port map( a => n5976, b => n5977, outb => 
                           mult_125_G3_FS_1_P_0_5_1_port);
   mult_125_G3_FS_1_U3_C_0_5_0 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_5_0_port, b => 
                           mult_125_G3_FS_1_C_1_5_0_port, outb => 
                           multiplier_sigs_2_22_port);
   mult_125_G3_FS_1_U3_B_0_5_0 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_5_0_port, b => 
                           mult_125_G3_FS_1_TEMP_P_0_5_0_port, outb => n5975);
   mult_125_G3_FS_1_U2_0_5_0 : nand2 port map( a => mult_125_G3_A1_20_port, b 
                           => mult_125_G3_A2_20_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_5_0_port);
   mult_125_G3_FS_1_U1_0_5_0 : nand2 port map( a => n5973, b => n5974, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_5_0_port);
   mult_125_G3_FS_1_U6_0_4_3 : oai12 port map( b => n5971, c => n5972, a => 
                           mult_125_G3_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G3_FS_1_C_1_4_3_port);
   mult_125_G3_FS_1_U5_0_4_3 : oai12 port map( b => n5969, c => n5970, a => 
                           mult_125_G3_FS_1_G_n_int_0_4_3_port, outb => 
                           mult_125_G3_FS_1_G_1_1_0_port);
   mult_125_G3_FS_1_U4_0_4_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_4_2_port, b => 
                           mult_125_G3_FS_1_P_0_4_3_port, outb => n6027);
   mult_125_G3_FS_1_U3_C_0_4_3 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_4_3_port, b => 
                           mult_125_G3_FS_1_C_1_4_3_port, outb => 
                           multiplier_sigs_2_21_port);
   mult_125_G3_FS_1_U3_B_0_4_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_4_3_port, b => 
                           mult_125_G3_FS_1_P_0_4_3_port, outb => n5968);
   mult_125_G3_FS_1_U2_0_4_3 : nand2 port map( a => mult_125_G3_A1_19_port, b 
                           => mult_125_G3_A2_19_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_4_3_port);
   mult_125_G3_FS_1_U1_0_4_3 : nand2 port map( a => n5966, b => n5967, outb => 
                           mult_125_G3_FS_1_P_0_4_3_port);
   mult_125_G3_FS_1_U6_0_4_2 : oai12 port map( b => n5964, c => n5965, a => 
                           mult_125_G3_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G3_FS_1_C_1_4_2_port);
   mult_125_G3_FS_1_U5_0_4_2 : oai12 port map( b => n5963, c => n5972, a => 
                           mult_125_G3_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_4_2_port);
   mult_125_G3_FS_1_U4_0_4_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_4_1_port, b => 
                           mult_125_G3_FS_1_P_0_4_2_port, outb => n5962);
   mult_125_G3_FS_1_U3_C_0_4_2 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_4_2_port, b => 
                           mult_125_G3_FS_1_C_1_4_2_port, outb => 
                           multiplier_sigs_2_20_port);
   mult_125_G3_FS_1_U3_B_0_4_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_4_2_port, b => 
                           mult_125_G3_FS_1_P_0_4_2_port, outb => n5961);
   mult_125_G3_FS_1_U2_0_4_2 : nand2 port map( a => mult_125_G3_A1_18_port, b 
                           => mult_125_G3_A2_18_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_4_2_port);
   mult_125_G3_FS_1_U1_0_4_2 : nand2 port map( a => n5959, b => n5960, outb => 
                           mult_125_G3_FS_1_P_0_4_2_port);
   mult_125_G3_FS_1_U6_0_4_1 : oai12 port map( b => n6026, c => n5958, a => 
                           mult_125_G3_FS_1_G_n_int_0_4_0_port, outb => 
                           mult_125_G3_FS_1_C_1_4_1_port);
   mult_125_G3_FS_1_U5_0_4_1 : oai12 port map( b => 
                           mult_125_G3_FS_1_G_n_int_0_4_0_port, c => n5965, a 
                           => mult_125_G3_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_4_1_port);
   mult_125_G3_FS_1_U4_0_4_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_TEMP_P_0_4_0_port, b => 
                           mult_125_G3_FS_1_P_0_4_1_port, outb => n5957);
   mult_125_G3_FS_1_U3_C_0_4_1 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_4_1_port, b => 
                           mult_125_G3_FS_1_C_1_4_1_port, outb => 
                           multiplier_sigs_2_19_port);
   mult_125_G3_FS_1_U3_B_0_4_1 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_4_1_port, b => 
                           mult_125_G3_FS_1_P_0_4_1_port, outb => n5956);
   mult_125_G3_FS_1_U2_0_4_1 : nand2 port map( a => mult_125_G3_A1_17_port, b 
                           => mult_125_G3_A2_17_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_4_1_port);
   mult_125_G3_FS_1_U1_0_4_1 : nand2 port map( a => n5954, b => n5955, outb => 
                           mult_125_G3_FS_1_P_0_4_1_port);
   mult_125_G3_FS_1_U3_C_0_4_0 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_4_0_port, b => 
                           mult_125_G3_FS_1_C_1_4_0_port, outb => 
                           multiplier_sigs_2_18_port);
   mult_125_G3_FS_1_U3_B_0_4_0 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_4_0_port, b => 
                           mult_125_G3_FS_1_TEMP_P_0_4_0_port, outb => n5953);
   mult_125_G3_FS_1_U2_0_4_0 : nand2 port map( a => mult_125_G3_A1_16_port, b 
                           => mult_125_G3_A2_16_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_4_0_port);
   mult_125_G3_FS_1_U1_0_4_0 : nand2 port map( a => n5951, b => n5952, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_4_0_port);
   mult_125_G3_FS_1_U5_0_3_3 : oai12 port map( b => n5949, c => n5950, a => 
                           mult_125_G3_FS_1_G_n_int_0_3_3_port, outb => 
                           mult_125_G3_FS_1_G_1_0_3_port);
   mult_125_G3_FS_1_U3_C_0_3_3 : xor2 port map( a => 
                           mult_125_G3_FS_1_PG_int_0_3_3_port, b => 
                           mult_125_G3_FS_1_C_1_3_3_port, outb => 
                           multiplier_sigs_2_17_port);
   mult_125_G3_FS_1_U3_B_0_3_3 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_3_3_port, b => 
                           mult_125_G3_FS_1_P_0_3_3_port, outb => n5948);
   mult_125_G3_FS_1_U2_0_3_3 : nand2 port map( a => mult_125_G3_A1_15_port, b 
                           => mult_125_G3_A2_15_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_3_3_port);
   mult_125_G3_FS_1_U1_0_3_3 : nand2 port map( a => n5946, b => n5947, outb => 
                           mult_125_G3_FS_1_P_0_3_3_port);
   mult_125_G3_FS_1_U3_B_0_3_2 : nand2 port map( a => 
                           mult_125_G3_FS_1_G_n_int_0_3_2_port, b => 
                           mult_125_G3_FS_1_P_0_3_2_port, outb => n5945);
   mult_125_G3_FS_1_U2_0_3_2 : nand2 port map( a => mult_125_G3_A1_14_port, b 
                           => mult_125_G3_A2_14_port, outb => 
                           mult_125_G3_FS_1_G_n_int_0_3_2_port);
   mult_125_G3_FS_1_U1_0_3_2 : nand2 port map( a => n5943, b => n5944, outb => 
                           mult_125_G3_FS_1_P_0_3_2_port);
   mult_125_G3_AN1_15 : inv port map( inb => coefficient_mem_array_2_15_port, 
                           outb => mult_125_G3_A_not_15_port);
   mult_125_G3_AN1_14 : inv port map( inb => coefficient_mem_array_2_14_port, 
                           outb => mult_125_G3_A_not_14_port);
   mult_125_G3_AN1_13 : inv port map( inb => coefficient_mem_array_2_13_port, 
                           outb => mult_125_G3_A_not_13_port);
   mult_125_G3_AN1_12 : inv port map( inb => coefficient_mem_array_2_12_port, 
                           outb => mult_125_G3_A_not_12_port);
   mult_125_G3_AN1_11 : inv port map( inb => coefficient_mem_array_2_11_port, 
                           outb => mult_125_G3_A_not_11_port);
   mult_125_G3_AN1_10 : inv port map( inb => coefficient_mem_array_2_10_port, 
                           outb => mult_125_G3_A_not_10_port);
   mult_125_G3_AN1_9 : inv port map( inb => coefficient_mem_array_2_9_port, 
                           outb => mult_125_G3_A_not_9_port);
   mult_125_G3_AN1_8 : inv port map( inb => coefficient_mem_array_2_8_port, 
                           outb => mult_125_G3_A_not_8_port);
   mult_125_G3_AN1_7 : inv port map( inb => coefficient_mem_array_2_7_port, 
                           outb => mult_125_G3_A_not_7_port);
   mult_125_G3_AN1_6 : inv port map( inb => coefficient_mem_array_2_6_port, 
                           outb => mult_125_G3_A_not_6_port);
   mult_125_G3_AN1_5 : inv port map( inb => coefficient_mem_array_2_5_port, 
                           outb => mult_125_G3_A_not_5_port);
   mult_125_G3_AN1_4 : inv port map( inb => coefficient_mem_array_2_4_port, 
                           outb => mult_125_G3_A_not_4_port);
   mult_125_G3_AN1_3 : inv port map( inb => coefficient_mem_array_2_3_port, 
                           outb => mult_125_G3_A_not_3_port);
   mult_125_G3_AN1_2 : inv port map( inb => coefficient_mem_array_2_2_port, 
                           outb => mult_125_G3_A_not_2_port);
   mult_125_G3_AN1_1 : inv port map( inb => coefficient_mem_array_2_1_port, 
                           outb => mult_125_G3_A_not_1_port);
   mult_125_G3_AN1_0 : inv port map( inb => coefficient_mem_array_2_0_port, 
                           outb => mult_125_G3_A_not_0_port);
   mult_125_G3_AN1_15_0 : inv port map( inb => input_sample_mem_15_port, outb 
                           => mult_125_G3_B_not_15_port);
   mult_125_G3_AN1_14_0 : inv port map( inb => input_sample_mem_14_port, outb 
                           => mult_125_G3_B_not_14_port);
   mult_125_G3_AN1_13_0 : inv port map( inb => input_sample_mem_13_port, outb 
                           => mult_125_G3_B_not_13_port);
   mult_125_G3_AN1_12_0 : inv port map( inb => input_sample_mem_12_port, outb 
                           => mult_125_G3_B_not_12_port);
   mult_125_G3_AN1_11_0 : inv port map( inb => input_sample_mem_11_port, outb 
                           => mult_125_G3_B_not_11_port);
   mult_125_G3_AN1_10_0 : inv port map( inb => input_sample_mem_10_port, outb 
                           => mult_125_G3_B_not_10_port);
   mult_125_G3_AN1_9_0 : inv port map( inb => input_sample_mem_9_port, outb => 
                           mult_125_G3_B_not_9_port);
   mult_125_G3_AN1_8_0 : inv port map( inb => input_sample_mem_8_port, outb => 
                           mult_125_G3_B_not_8_port);
   mult_125_G3_AN1_7_0 : inv port map( inb => input_sample_mem_7_port, outb => 
                           mult_125_G3_B_not_7_port);
   mult_125_G3_AN1_6_0 : inv port map( inb => input_sample_mem_6_port, outb => 
                           mult_125_G3_B_not_6_port);
   mult_125_G3_AN1_5_0 : inv port map( inb => input_sample_mem_5_port, outb => 
                           mult_125_G3_B_not_5_port);
   mult_125_G3_AN1_4_0 : inv port map( inb => input_sample_mem_4_port, outb => 
                           mult_125_G3_B_not_4_port);
   mult_125_G3_AN1_3_0 : inv port map( inb => input_sample_mem_3_port, outb => 
                           mult_125_G3_B_not_3_port);
   mult_125_G3_AN1_2_0 : inv port map( inb => input_sample_mem_2_port, outb => 
                           mult_125_G3_B_not_2_port);
   mult_125_G3_AN1_1_0 : inv port map( inb => input_sample_mem_1_port, outb => 
                           mult_125_G3_B_not_1_port);
   mult_125_G3_AN1_0_0 : inv port map( inb => input_sample_mem_0_port, outb => 
                           mult_125_G3_B_not_0_port);
   mult_125_G3_AN1_15_15 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_15_15_port);
   mult_125_G3_AN3_15_14 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_14_port, outb => 
                           mult_125_G3_ab_15_14_port);
   mult_125_G3_AN3_15_13 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_13_port, outb => 
                           mult_125_G3_ab_15_13_port);
   mult_125_G3_AN3_15_12 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_12_port, outb => 
                           mult_125_G3_ab_15_12_port);
   mult_125_G3_AN3_15_11 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_11_port, outb => 
                           mult_125_G3_ab_15_11_port);
   mult_125_G3_AN3_15_10 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_10_port, outb => 
                           mult_125_G3_ab_15_10_port);
   mult_125_G3_AN3_15_9 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_9_port, outb => 
                           mult_125_G3_ab_15_9_port);
   mult_125_G3_AN3_15_8 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_8_port, outb => 
                           mult_125_G3_ab_15_8_port);
   mult_125_G3_AN3_15_7 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_7_port, outb => 
                           mult_125_G3_ab_15_7_port);
   mult_125_G3_AN3_15_6 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_6_port, outb => 
                           mult_125_G3_ab_15_6_port);
   mult_125_G3_AN3_15_5 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_5_port, outb => 
                           mult_125_G3_ab_15_5_port);
   mult_125_G3_AN3_15_4 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_4_port, outb => 
                           mult_125_G3_ab_15_4_port);
   mult_125_G3_AN3_15_3 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_3_port, outb => 
                           mult_125_G3_ab_15_3_port);
   mult_125_G3_AN3_15_2 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_2_port, outb => 
                           mult_125_G3_ab_15_2_port);
   mult_125_G3_AN3_15_1 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_1_port, outb => 
                           mult_125_G3_ab_15_1_port);
   mult_125_G3_AN3_15_0 : nor2 port map( a => mult_125_G3_A_not_15_port, b => 
                           mult_125_G3_B_notx_0_port, outb => 
                           mult_125_G3_ab_15_0_port);
   mult_125_G3_AN2_14_15 : nor2 port map( a => mult_125_G3_A_notx_14_port, b =>
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_14_15_port);
   mult_125_G3_AN1_14_14 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_14_14_port);
   mult_125_G3_AN1_14_13 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_14_13_port);
   mult_125_G3_AN1_14_12 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_14_12_port);
   mult_125_G3_AN1_14_11 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_14_11_port);
   mult_125_G3_AN1_14_10 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_14_10_port);
   mult_125_G3_AN1_14_9 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_14_9_port);
   mult_125_G3_AN1_14_8 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_14_8_port);
   mult_125_G3_AN1_14_7 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_14_7_port);
   mult_125_G3_AN1_14_6 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_14_6_port);
   mult_125_G3_AN1_14_5 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_14_5_port);
   mult_125_G3_AN1_14_4 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_14_4_port);
   mult_125_G3_AN1_14_3 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_14_3_port);
   mult_125_G3_AN1_14_2 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_14_2_port);
   mult_125_G3_AN1_14_1 : nor2 port map( a => mult_125_G3_A_not_14_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_14_1_port);
   mult_125_G3_AN1_14_0_0 : nor2 port map( a => mult_125_G3_A_not_14_port, b =>
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_14_0_port);
   mult_125_G3_AN2_13_15 : nor2 port map( a => mult_125_G3_A_notx_13_port, b =>
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_13_15_port);
   mult_125_G3_AN1_13_14 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_13_14_port);
   mult_125_G3_AN1_13_13 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_13_13_port);
   mult_125_G3_AN1_13_12 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_13_12_port);
   mult_125_G3_AN1_13_11 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_13_11_port);
   mult_125_G3_AN1_13_10 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_13_10_port);
   mult_125_G3_AN1_13_9 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_13_9_port);
   mult_125_G3_AN1_13_8 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_13_8_port);
   mult_125_G3_AN1_13_7 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_13_7_port);
   mult_125_G3_AN1_13_6 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_13_6_port);
   mult_125_G3_AN1_13_5 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_13_5_port);
   mult_125_G3_AN1_13_4 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_13_4_port);
   mult_125_G3_AN1_13_3 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_13_3_port);
   mult_125_G3_AN1_13_2 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_13_2_port);
   mult_125_G3_AN1_13_1 : nor2 port map( a => mult_125_G3_A_not_13_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_13_1_port);
   mult_125_G3_AN1_13_0_0 : nor2 port map( a => mult_125_G3_A_not_13_port, b =>
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_13_0_port);
   mult_125_G3_AN2_12_15 : nor2 port map( a => mult_125_G3_A_notx_12_port, b =>
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_12_15_port);
   mult_125_G3_AN1_12_14 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_12_14_port);
   mult_125_G3_AN1_12_13 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_12_13_port);
   mult_125_G3_AN1_12_12 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_12_12_port);
   mult_125_G3_AN1_12_11 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_12_11_port);
   mult_125_G3_AN1_12_10 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_12_10_port);
   mult_125_G3_AN1_12_9 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_12_9_port);
   mult_125_G3_AN1_12_8 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_12_8_port);
   mult_125_G3_AN1_12_7 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_12_7_port);
   mult_125_G3_AN1_12_6 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_12_6_port);
   mult_125_G3_AN1_12_5 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_12_5_port);
   mult_125_G3_AN1_12_4 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_12_4_port);
   mult_125_G3_AN1_12_3 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_12_3_port);
   mult_125_G3_AN1_12_2 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_12_2_port);
   mult_125_G3_AN1_12_1 : nor2 port map( a => mult_125_G3_A_not_12_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_12_1_port);
   mult_125_G3_AN1_12_0_0 : nor2 port map( a => mult_125_G3_A_not_12_port, b =>
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_12_0_port);
   mult_125_G3_AN2_11_15 : nor2 port map( a => mult_125_G3_A_notx_11_port, b =>
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_11_15_port);
   mult_125_G3_AN1_11_14 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_11_14_port);
   mult_125_G3_AN1_11_13 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_11_13_port);
   mult_125_G3_AN1_11_12 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_11_12_port);
   mult_125_G3_AN1_11_11 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_11_11_port);
   mult_125_G3_AN1_11_10 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_11_10_port);
   mult_125_G3_AN1_11_9 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_11_9_port);
   mult_125_G3_AN1_11_8 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_11_8_port);
   mult_125_G3_AN1_11_7 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_11_7_port);
   mult_125_G3_AN1_11_6 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_11_6_port);
   mult_125_G3_AN1_11_5 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_11_5_port);
   mult_125_G3_AN1_11_4 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_11_4_port);
   mult_125_G3_AN1_11_3 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_11_3_port);
   mult_125_G3_AN1_11_2 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_11_2_port);
   mult_125_G3_AN1_11_1 : nor2 port map( a => mult_125_G3_A_not_11_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_11_1_port);
   mult_125_G3_AN1_11_0_0 : nor2 port map( a => mult_125_G3_A_not_11_port, b =>
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_11_0_port);
   mult_125_G3_AN2_10_15 : nor2 port map( a => mult_125_G3_A_notx_10_port, b =>
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_10_15_port);
   mult_125_G3_AN1_10_14 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_10_14_port);
   mult_125_G3_AN1_10_13 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_10_13_port);
   mult_125_G3_AN1_10_12 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_10_12_port);
   mult_125_G3_AN1_10_11 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_10_11_port);
   mult_125_G3_AN1_10_10 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_10_10_port);
   mult_125_G3_AN1_10_9 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_10_9_port);
   mult_125_G3_AN1_10_8 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_10_8_port);
   mult_125_G3_AN1_10_7 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_10_7_port);
   mult_125_G3_AN1_10_6 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_10_6_port);
   mult_125_G3_AN1_10_5 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_10_5_port);
   mult_125_G3_AN1_10_4 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_10_4_port);
   mult_125_G3_AN1_10_3 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_10_3_port);
   mult_125_G3_AN1_10_2 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_10_2_port);
   mult_125_G3_AN1_10_1 : nor2 port map( a => mult_125_G3_A_not_10_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_10_1_port);
   mult_125_G3_AN1_10_0_0 : nor2 port map( a => mult_125_G3_A_not_10_port, b =>
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_10_0_port);
   mult_125_G3_AN2_9_15 : nor2 port map( a => mult_125_G3_A_notx_9_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_9_15_port);
   mult_125_G3_AN1_9_14 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_9_14_port);
   mult_125_G3_AN1_9_13 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_9_13_port);
   mult_125_G3_AN1_9_12 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_9_12_port);
   mult_125_G3_AN1_9_11 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_9_11_port);
   mult_125_G3_AN1_9_10 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_9_10_port);
   mult_125_G3_AN1_9_9 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_9_9_port);
   mult_125_G3_AN1_9_8 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_9_8_port);
   mult_125_G3_AN1_9_7 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_9_7_port);
   mult_125_G3_AN1_9_6 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_9_6_port);
   mult_125_G3_AN1_9_5 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_9_5_port);
   mult_125_G3_AN1_9_4 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_9_4_port);
   mult_125_G3_AN1_9_3 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_9_3_port);
   mult_125_G3_AN1_9_2 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_9_2_port);
   mult_125_G3_AN1_9_1 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_9_1_port);
   mult_125_G3_AN1_9_0_0 : nor2 port map( a => mult_125_G3_A_not_9_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_9_0_port);
   mult_125_G3_AN2_8_15 : nor2 port map( a => mult_125_G3_A_notx_8_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_8_15_port);
   mult_125_G3_AN1_8_14 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_8_14_port);
   mult_125_G3_AN1_8_13 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_8_13_port);
   mult_125_G3_AN1_8_12 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_8_12_port);
   mult_125_G3_AN1_8_11 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_8_11_port);
   mult_125_G3_AN1_8_10 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_8_10_port);
   mult_125_G3_AN1_8_9 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_8_9_port);
   mult_125_G3_AN1_8_8 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_8_8_port);
   mult_125_G3_AN1_8_7 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_8_7_port);
   mult_125_G3_AN1_8_6 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_8_6_port);
   mult_125_G3_AN1_8_5 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_8_5_port);
   mult_125_G3_AN1_8_4 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_8_4_port);
   mult_125_G3_AN1_8_3 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_8_3_port);
   mult_125_G3_AN1_8_2 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_8_2_port);
   mult_125_G3_AN1_8_1 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_8_1_port);
   mult_125_G3_AN1_8_0_0 : nor2 port map( a => mult_125_G3_A_not_8_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_8_0_port);
   mult_125_G3_AN2_7_15 : nor2 port map( a => mult_125_G3_A_notx_7_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_7_15_port);
   mult_125_G3_AN1_7_14 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_7_14_port);
   mult_125_G3_AN1_7_13 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_7_13_port);
   mult_125_G3_AN1_7_12 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_7_12_port);
   mult_125_G3_AN1_7_11 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_7_11_port);
   mult_125_G3_AN1_7_10 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_7_10_port);
   mult_125_G3_AN1_7_9 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_7_9_port);
   mult_125_G3_AN1_7_8 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_7_8_port);
   mult_125_G3_AN1_7_7 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_7_7_port);
   mult_125_G3_AN1_7_6 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_7_6_port);
   mult_125_G3_AN1_7_5 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_7_5_port);
   mult_125_G3_AN1_7_4 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_7_4_port);
   mult_125_G3_AN1_7_3 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_7_3_port);
   mult_125_G3_AN1_7_2 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_7_2_port);
   mult_125_G3_AN1_7_1 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_7_1_port);
   mult_125_G3_AN1_7_0_0 : nor2 port map( a => mult_125_G3_A_not_7_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_7_0_port);
   mult_125_G3_AN2_6_15 : nor2 port map( a => mult_125_G3_A_notx_6_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_6_15_port);
   mult_125_G3_AN1_6_14 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_6_14_port);
   mult_125_G3_AN1_6_13 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_6_13_port);
   mult_125_G3_AN1_6_12 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_6_12_port);
   mult_125_G3_AN1_6_11 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_6_11_port);
   mult_125_G3_AN1_6_10 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_6_10_port);
   mult_125_G3_AN1_6_9 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_6_9_port);
   mult_125_G3_AN1_6_8 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_6_8_port);
   mult_125_G3_AN1_6_7 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_6_7_port);
   mult_125_G3_AN1_6_6 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_6_6_port);
   mult_125_G3_AN1_6_5 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_6_5_port);
   mult_125_G3_AN1_6_4 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_6_4_port);
   mult_125_G3_AN1_6_3 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_6_3_port);
   mult_125_G3_AN1_6_2 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_6_2_port);
   mult_125_G3_AN1_6_1 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_6_1_port);
   mult_125_G3_AN1_6_0_0 : nor2 port map( a => mult_125_G3_A_not_6_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_6_0_port);
   mult_125_G3_AN2_5_15 : nor2 port map( a => mult_125_G3_A_notx_5_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_5_15_port);
   mult_125_G3_AN1_5_14 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_5_14_port);
   mult_125_G3_AN1_5_13 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_5_13_port);
   mult_125_G3_AN1_5_12 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_5_12_port);
   mult_125_G3_AN1_5_11 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_5_11_port);
   mult_125_G3_AN1_5_10 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_5_10_port);
   mult_125_G3_AN1_5_9 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_5_9_port);
   mult_125_G3_AN1_5_8 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_5_8_port);
   mult_125_G3_AN1_5_7 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_5_7_port);
   mult_125_G3_AN1_5_6 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_5_6_port);
   mult_125_G3_AN1_5_5 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_5_5_port);
   mult_125_G3_AN1_5_4 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_5_4_port);
   mult_125_G3_AN1_5_3 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_5_3_port);
   mult_125_G3_AN1_5_2 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_5_2_port);
   mult_125_G3_AN1_5_1 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_5_1_port);
   mult_125_G3_AN1_5_0_0 : nor2 port map( a => mult_125_G3_A_not_5_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_5_0_port);
   mult_125_G3_AN2_4_15 : nor2 port map( a => mult_125_G3_A_notx_4_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_4_15_port);
   mult_125_G3_AN1_4_14 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_4_14_port);
   mult_125_G3_AN1_4_13 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_4_13_port);
   mult_125_G3_AN1_4_12 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_4_12_port);
   mult_125_G3_AN1_4_11 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_4_11_port);
   mult_125_G3_AN1_4_10 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_4_10_port);
   mult_125_G3_AN1_4_9 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_4_9_port);
   mult_125_G3_AN1_4_8 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_4_8_port);
   mult_125_G3_AN1_4_7 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_4_7_port);
   mult_125_G3_AN1_4_6 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_4_6_port);
   mult_125_G3_AN1_4_5 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_4_5_port);
   mult_125_G3_AN1_4_4 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_4_4_port);
   mult_125_G3_AN1_4_3 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_4_3_port);
   mult_125_G3_AN1_4_2 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_4_2_port);
   mult_125_G3_AN1_4_1 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_4_1_port);
   mult_125_G3_AN1_4_0_0 : nor2 port map( a => mult_125_G3_A_not_4_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_4_0_port);
   mult_125_G3_AN2_3_15 : nor2 port map( a => mult_125_G3_A_notx_3_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_3_15_port);
   mult_125_G3_AN1_3_14 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_3_14_port);
   mult_125_G3_AN1_3_13 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_3_13_port);
   mult_125_G3_AN1_3_12 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_3_12_port);
   mult_125_G3_AN1_3_11 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_3_11_port);
   mult_125_G3_AN1_3_10 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_3_10_port);
   mult_125_G3_AN1_3_9 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_3_9_port);
   mult_125_G3_AN1_3_8 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_3_8_port);
   mult_125_G3_AN1_3_7 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_3_7_port);
   mult_125_G3_AN1_3_6 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_3_6_port);
   mult_125_G3_AN1_3_5 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_3_5_port);
   mult_125_G3_AN1_3_4 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_3_4_port);
   mult_125_G3_AN1_3_3 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_3_3_port);
   mult_125_G3_AN1_3_2 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_3_2_port);
   mult_125_G3_AN1_3_1 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_3_1_port);
   mult_125_G3_AN1_3_0_0 : nor2 port map( a => mult_125_G3_A_not_3_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_3_0_port);
   mult_125_G3_AN2_2_15 : nor2 port map( a => mult_125_G3_A_notx_2_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_2_15_port);
   mult_125_G3_AN1_2_14 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_2_14_port);
   mult_125_G3_AN1_2_13 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_2_13_port);
   mult_125_G3_AN1_2_12 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_2_12_port);
   mult_125_G3_AN1_2_11 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_2_11_port);
   mult_125_G3_AN1_2_10 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_2_10_port);
   mult_125_G3_AN1_2_9 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_2_9_port);
   mult_125_G3_AN1_2_8 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_2_8_port);
   mult_125_G3_AN1_2_7 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_2_7_port);
   mult_125_G3_AN1_2_6 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_2_6_port);
   mult_125_G3_AN1_2_5 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_2_5_port);
   mult_125_G3_AN1_2_4 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_2_4_port);
   mult_125_G3_AN1_2_3 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_2_3_port);
   mult_125_G3_AN1_2_2 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_2_2_port);
   mult_125_G3_AN1_2_1 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_2_1_port);
   mult_125_G3_AN1_2_0_0 : nor2 port map( a => mult_125_G3_A_not_2_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_2_0_port);
   mult_125_G3_AN2_1_15 : nor2 port map( a => mult_125_G3_A_notx_1_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_1_15_port);
   mult_125_G3_AN1_1_14 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_1_14_port);
   mult_125_G3_AN1_1_13 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_1_13_port);
   mult_125_G3_AN1_1_12 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_1_12_port);
   mult_125_G3_AN1_1_11 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_1_11_port);
   mult_125_G3_AN1_1_10 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_1_10_port);
   mult_125_G3_AN1_1_9 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_1_9_port);
   mult_125_G3_AN1_1_8 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_1_8_port);
   mult_125_G3_AN1_1_7 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_1_7_port);
   mult_125_G3_AN1_1_6 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_1_6_port);
   mult_125_G3_AN1_1_5 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_1_5_port);
   mult_125_G3_AN1_1_4 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_1_4_port);
   mult_125_G3_AN1_1_3 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_1_3_port);
   mult_125_G3_AN1_1_2 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_1_2_port);
   mult_125_G3_AN1_1_1 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_1_1_port);
   mult_125_G3_AN1_1_0_0 : nor2 port map( a => mult_125_G3_A_not_1_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_ab_1_0_port);
   mult_125_G3_AN2_0_15 : nor2 port map( a => mult_125_G3_A_notx_0_port, b => 
                           mult_125_G3_B_not_15_port, outb => 
                           mult_125_G3_ab_0_15_port);
   mult_125_G3_AN1_0_14 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_ab_0_14_port);
   mult_125_G3_AN1_0_13 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_ab_0_13_port);
   mult_125_G3_AN1_0_12 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_ab_0_12_port);
   mult_125_G3_AN1_0_11 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_ab_0_11_port);
   mult_125_G3_AN1_0_10 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_ab_0_10_port);
   mult_125_G3_AN1_0_9 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_ab_0_9_port);
   mult_125_G3_AN1_0_8 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_ab_0_8_port);
   mult_125_G3_AN1_0_7 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_ab_0_7_port);
   mult_125_G3_AN1_0_6 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_ab_0_6_port);
   mult_125_G3_AN1_0_5 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_ab_0_5_port);
   mult_125_G3_AN1_0_4 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_ab_0_4_port);
   mult_125_G3_AN1_0_3 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_ab_0_3_port);
   mult_125_G3_AN1_0_2 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_ab_0_2_port);
   mult_125_G3_AN1_0_1 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_ab_0_1_port);
   mult_125_G3_AN1_0_0_0 : nor2 port map( a => mult_125_G3_A_not_0_port, b => 
                           mult_125_G3_B_not_0_port, outb => 
                           multiplier_sigs_2_0_port);
   mult_125_G2_FS_1_U6_1_1_3 : oai12 port map( b => n5907, c => n5908, a => 
                           n5909, outb => mult_125_G2_FS_1_C_1_7_0_port);
   mult_125_G2_FS_1_U6_1_1_2 : oai12 port map( b => n5904, c => n5905, a => 
                           n5906, outb => mult_125_G2_FS_1_C_1_6_0_port);
   mult_125_G2_FS_1_U6_1_1_1 : oai12 port map( b => n5901, c => n5902, a => 
                           n5903, outb => mult_125_G2_FS_1_C_1_5_0_port);
   mult_125_G2_FS_1_U6_0_7_1 : oai12 port map( b => n5898, c => n5899, a => 
                           mult_125_G2_FS_1_G_n_int_0_7_0_port, outb => 
                           mult_125_G2_FS_1_C_1_7_1_port);
   mult_125_G2_FS_1_U3_C_0_7_1 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_7_1_port, b => 
                           mult_125_G2_FS_1_C_1_7_1_port, outb => 
                           multiplier_sigs_1_31_port);
   mult_125_G2_FS_1_U3_B_0_7_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_7_1_port, b => 
                           mult_125_G2_FS_1_P_0_7_1_port, outb => n5897);
   mult_125_G2_FS_1_U2_0_7_1 : nand2 port map( a => mult_125_G2_A1_29_port, b 
                           => mult_125_G2_A2_29_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_7_1_port);
   mult_125_G2_FS_1_U1_0_7_1 : nand2 port map( a => n5895, b => n5896, outb => 
                           mult_125_G2_FS_1_P_0_7_1_port);
   mult_125_G2_FS_1_U3_C_0_7_0 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_7_0_port, b => 
                           mult_125_G2_FS_1_C_1_7_0_port, outb => 
                           multiplier_sigs_1_30_port);
   mult_125_G2_FS_1_U3_B_0_7_0 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_7_0_port, b => 
                           mult_125_G2_FS_1_TEMP_P_0_7_0_port, outb => n5894);
   mult_125_G2_FS_1_U2_0_7_0 : nand2 port map( a => mult_125_G2_A1_28_port, b 
                           => mult_125_G2_A2_28_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_7_0_port);
   mult_125_G2_FS_1_U1_0_7_0 : nand2 port map( a => n5892, b => n5893, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_7_0_port);
   mult_125_G2_FS_1_U6_0_6_3 : oai12 port map( b => n5890, c => n5891, a => 
                           mult_125_G2_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G2_FS_1_C_1_6_3_port);
   mult_125_G2_FS_1_U5_0_6_3 : oai12 port map( b => n5888, c => n5889, a => 
                           mult_125_G2_FS_1_G_n_int_0_6_3_port, outb => 
                           mult_125_G2_FS_1_G_1_1_2_port);
   mult_125_G2_FS_1_U4_0_6_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_6_2_port, b => 
                           mult_125_G2_FS_1_P_0_6_3_port, outb => n5908);
   mult_125_G2_FS_1_U3_C_0_6_3 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_6_3_port, b => 
                           mult_125_G2_FS_1_C_1_6_3_port, outb => 
                           multiplier_sigs_1_29_port);
   mult_125_G2_FS_1_U3_B_0_6_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_6_3_port, b => 
                           mult_125_G2_FS_1_P_0_6_3_port, outb => n5887);
   mult_125_G2_FS_1_U2_0_6_3 : nand2 port map( a => mult_125_G2_A1_27_port, b 
                           => mult_125_G2_A2_27_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_6_3_port);
   mult_125_G2_FS_1_U1_0_6_3 : nand2 port map( a => n5885, b => n5886, outb => 
                           mult_125_G2_FS_1_P_0_6_3_port);
   mult_125_G2_FS_1_U6_0_6_2 : oai12 port map( b => n5883, c => n5884, a => 
                           mult_125_G2_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G2_FS_1_C_1_6_2_port);
   mult_125_G2_FS_1_U5_0_6_2 : oai12 port map( b => n5882, c => n5891, a => 
                           mult_125_G2_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_6_2_port);
   mult_125_G2_FS_1_U4_0_6_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_6_1_port, b => 
                           mult_125_G2_FS_1_P_0_6_2_port, outb => n5881);
   mult_125_G2_FS_1_U3_C_0_6_2 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_6_2_port, b => 
                           mult_125_G2_FS_1_C_1_6_2_port, outb => 
                           multiplier_sigs_1_28_port);
   mult_125_G2_FS_1_U3_B_0_6_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_6_2_port, b => 
                           mult_125_G2_FS_1_P_0_6_2_port, outb => n5880);
   mult_125_G2_FS_1_U2_0_6_2 : nand2 port map( a => mult_125_G2_A1_26_port, b 
                           => mult_125_G2_A2_26_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_6_2_port);
   mult_125_G2_FS_1_U1_0_6_2 : nand2 port map( a => n5878, b => n5879, outb => 
                           mult_125_G2_FS_1_P_0_6_2_port);
   mult_125_G2_FS_1_U6_0_6_1 : oai12 port map( b => n5907, c => n5877, a => 
                           mult_125_G2_FS_1_G_n_int_0_6_0_port, outb => 
                           mult_125_G2_FS_1_C_1_6_1_port);
   mult_125_G2_FS_1_U5_0_6_1 : oai12 port map( b => 
                           mult_125_G2_FS_1_G_n_int_0_6_0_port, c => n5884, a 
                           => mult_125_G2_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_6_1_port);
   mult_125_G2_FS_1_U4_0_6_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_6_0_port, b => 
                           mult_125_G2_FS_1_P_0_6_1_port, outb => n5876);
   mult_125_G2_FS_1_U3_C_0_6_1 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_6_1_port, b => 
                           mult_125_G2_FS_1_C_1_6_1_port, outb => 
                           multiplier_sigs_1_27_port);
   mult_125_G2_FS_1_U3_B_0_6_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_6_1_port, b => 
                           mult_125_G2_FS_1_P_0_6_1_port, outb => n5875);
   mult_125_G2_FS_1_U2_0_6_1 : nand2 port map( a => mult_125_G2_A1_25_port, b 
                           => mult_125_G2_A2_25_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_6_1_port);
   mult_125_G2_FS_1_U1_0_6_1 : nand2 port map( a => n5873, b => n5874, outb => 
                           mult_125_G2_FS_1_P_0_6_1_port);
   mult_125_G2_FS_1_U3_C_0_6_0 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_6_0_port, b => 
                           mult_125_G2_FS_1_C_1_6_0_port, outb => 
                           multiplier_sigs_1_26_port);
   mult_125_G2_FS_1_U3_B_0_6_0 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_6_0_port, b => 
                           mult_125_G2_FS_1_TEMP_P_0_6_0_port, outb => n5872);
   mult_125_G2_FS_1_U2_0_6_0 : nand2 port map( a => mult_125_G2_A1_24_port, b 
                           => mult_125_G2_A2_24_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_6_0_port);
   mult_125_G2_FS_1_U1_0_6_0 : nand2 port map( a => n5870, b => n5871, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_6_0_port);
   mult_125_G2_FS_1_U6_0_5_3 : oai12 port map( b => n5868, c => n5869, a => 
                           mult_125_G2_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G2_FS_1_C_1_5_3_port);
   mult_125_G2_FS_1_U5_0_5_3 : oai12 port map( b => n5866, c => n5867, a => 
                           mult_125_G2_FS_1_G_n_int_0_5_3_port, outb => 
                           mult_125_G2_FS_1_G_1_1_1_port);
   mult_125_G2_FS_1_U4_0_5_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_5_2_port, b => 
                           mult_125_G2_FS_1_P_0_5_3_port, outb => n5905);
   mult_125_G2_FS_1_U3_C_0_5_3 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_5_3_port, b => 
                           mult_125_G2_FS_1_C_1_5_3_port, outb => 
                           multiplier_sigs_1_25_port);
   mult_125_G2_FS_1_U3_B_0_5_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_5_3_port, b => 
                           mult_125_G2_FS_1_P_0_5_3_port, outb => n5865);
   mult_125_G2_FS_1_U2_0_5_3 : nand2 port map( a => mult_125_G2_A1_23_port, b 
                           => mult_125_G2_A2_23_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_5_3_port);
   mult_125_G2_FS_1_U1_0_5_3 : nand2 port map( a => n5863, b => n5864, outb => 
                           mult_125_G2_FS_1_P_0_5_3_port);
   mult_125_G2_FS_1_U6_0_5_2 : oai12 port map( b => n5861, c => n5862, a => 
                           mult_125_G2_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G2_FS_1_C_1_5_2_port);
   mult_125_G2_FS_1_U5_0_5_2 : oai12 port map( b => n5860, c => n5869, a => 
                           mult_125_G2_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_5_2_port);
   mult_125_G2_FS_1_U4_0_5_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_5_1_port, b => 
                           mult_125_G2_FS_1_P_0_5_2_port, outb => n5859);
   mult_125_G2_FS_1_U3_C_0_5_2 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_5_2_port, b => 
                           mult_125_G2_FS_1_C_1_5_2_port, outb => 
                           multiplier_sigs_1_24_port);
   mult_125_G2_FS_1_U3_B_0_5_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_5_2_port, b => 
                           mult_125_G2_FS_1_P_0_5_2_port, outb => n5858);
   mult_125_G2_FS_1_U2_0_5_2 : nand2 port map( a => mult_125_G2_A1_22_port, b 
                           => mult_125_G2_A2_22_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_5_2_port);
   mult_125_G2_FS_1_U1_0_5_2 : nand2 port map( a => n5856, b => n5857, outb => 
                           mult_125_G2_FS_1_P_0_5_2_port);
   mult_125_G2_FS_1_U6_0_5_1 : oai12 port map( b => n5904, c => n5855, a => 
                           mult_125_G2_FS_1_G_n_int_0_5_0_port, outb => 
                           mult_125_G2_FS_1_C_1_5_1_port);
   mult_125_G2_FS_1_U5_0_5_1 : oai12 port map( b => 
                           mult_125_G2_FS_1_G_n_int_0_5_0_port, c => n5862, a 
                           => mult_125_G2_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_5_1_port);
   mult_125_G2_FS_1_U4_0_5_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_5_0_port, b => 
                           mult_125_G2_FS_1_P_0_5_1_port, outb => n5854);
   mult_125_G2_FS_1_U3_C_0_5_1 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_5_1_port, b => 
                           mult_125_G2_FS_1_C_1_5_1_port, outb => 
                           multiplier_sigs_1_23_port);
   mult_125_G2_FS_1_U3_B_0_5_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_5_1_port, b => 
                           mult_125_G2_FS_1_P_0_5_1_port, outb => n5853);
   mult_125_G2_FS_1_U2_0_5_1 : nand2 port map( a => mult_125_G2_A1_21_port, b 
                           => mult_125_G2_A2_21_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_5_1_port);
   mult_125_G2_FS_1_U1_0_5_1 : nand2 port map( a => n5851, b => n5852, outb => 
                           mult_125_G2_FS_1_P_0_5_1_port);
   mult_125_G2_FS_1_U3_C_0_5_0 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_5_0_port, b => 
                           mult_125_G2_FS_1_C_1_5_0_port, outb => 
                           multiplier_sigs_1_22_port);
   mult_125_G2_FS_1_U3_B_0_5_0 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_5_0_port, b => 
                           mult_125_G2_FS_1_TEMP_P_0_5_0_port, outb => n5850);
   mult_125_G2_FS_1_U2_0_5_0 : nand2 port map( a => mult_125_G2_A1_20_port, b 
                           => mult_125_G2_A2_20_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_5_0_port);
   mult_125_G2_FS_1_U1_0_5_0 : nand2 port map( a => n5848, b => n5849, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_5_0_port);
   mult_125_G2_FS_1_U6_0_4_3 : oai12 port map( b => n5846, c => n5847, a => 
                           mult_125_G2_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G2_FS_1_C_1_4_3_port);
   mult_125_G2_FS_1_U5_0_4_3 : oai12 port map( b => n5844, c => n5845, a => 
                           mult_125_G2_FS_1_G_n_int_0_4_3_port, outb => 
                           mult_125_G2_FS_1_G_1_1_0_port);
   mult_125_G2_FS_1_U4_0_4_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_4_2_port, b => 
                           mult_125_G2_FS_1_P_0_4_3_port, outb => n5902);
   mult_125_G2_FS_1_U3_C_0_4_3 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_4_3_port, b => 
                           mult_125_G2_FS_1_C_1_4_3_port, outb => 
                           multiplier_sigs_1_21_port);
   mult_125_G2_FS_1_U3_B_0_4_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_4_3_port, b => 
                           mult_125_G2_FS_1_P_0_4_3_port, outb => n5843);
   mult_125_G2_FS_1_U2_0_4_3 : nand2 port map( a => mult_125_G2_A1_19_port, b 
                           => mult_125_G2_A2_19_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_4_3_port);
   mult_125_G2_FS_1_U1_0_4_3 : nand2 port map( a => n5841, b => n5842, outb => 
                           mult_125_G2_FS_1_P_0_4_3_port);
   mult_125_G2_FS_1_U6_0_4_2 : oai12 port map( b => n5839, c => n5840, a => 
                           mult_125_G2_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G2_FS_1_C_1_4_2_port);
   mult_125_G2_FS_1_U5_0_4_2 : oai12 port map( b => n5838, c => n5847, a => 
                           mult_125_G2_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_4_2_port);
   mult_125_G2_FS_1_U4_0_4_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_4_1_port, b => 
                           mult_125_G2_FS_1_P_0_4_2_port, outb => n5837);
   mult_125_G2_FS_1_U3_C_0_4_2 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_4_2_port, b => 
                           mult_125_G2_FS_1_C_1_4_2_port, outb => 
                           multiplier_sigs_1_20_port);
   mult_125_G2_FS_1_U3_B_0_4_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_4_2_port, b => 
                           mult_125_G2_FS_1_P_0_4_2_port, outb => n5836);
   mult_125_G2_FS_1_U2_0_4_2 : nand2 port map( a => mult_125_G2_A1_18_port, b 
                           => mult_125_G2_A2_18_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_4_2_port);
   mult_125_G2_FS_1_U1_0_4_2 : nand2 port map( a => n5834, b => n5835, outb => 
                           mult_125_G2_FS_1_P_0_4_2_port);
   mult_125_G2_FS_1_U6_0_4_1 : oai12 port map( b => n5901, c => n5833, a => 
                           mult_125_G2_FS_1_G_n_int_0_4_0_port, outb => 
                           mult_125_G2_FS_1_C_1_4_1_port);
   mult_125_G2_FS_1_U5_0_4_1 : oai12 port map( b => 
                           mult_125_G2_FS_1_G_n_int_0_4_0_port, c => n5840, a 
                           => mult_125_G2_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_4_1_port);
   mult_125_G2_FS_1_U4_0_4_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_TEMP_P_0_4_0_port, b => 
                           mult_125_G2_FS_1_P_0_4_1_port, outb => n5832);
   mult_125_G2_FS_1_U3_C_0_4_1 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_4_1_port, b => 
                           mult_125_G2_FS_1_C_1_4_1_port, outb => 
                           multiplier_sigs_1_19_port);
   mult_125_G2_FS_1_U3_B_0_4_1 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_4_1_port, b => 
                           mult_125_G2_FS_1_P_0_4_1_port, outb => n5831);
   mult_125_G2_FS_1_U2_0_4_1 : nand2 port map( a => mult_125_G2_A1_17_port, b 
                           => mult_125_G2_A2_17_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_4_1_port);
   mult_125_G2_FS_1_U1_0_4_1 : nand2 port map( a => n5829, b => n5830, outb => 
                           mult_125_G2_FS_1_P_0_4_1_port);
   mult_125_G2_FS_1_U3_C_0_4_0 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_4_0_port, b => 
                           mult_125_G2_FS_1_C_1_4_0_port, outb => 
                           multiplier_sigs_1_18_port);
   mult_125_G2_FS_1_U3_B_0_4_0 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_4_0_port, b => 
                           mult_125_G2_FS_1_TEMP_P_0_4_0_port, outb => n5828);
   mult_125_G2_FS_1_U2_0_4_0 : nand2 port map( a => mult_125_G2_A1_16_port, b 
                           => mult_125_G2_A2_16_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_4_0_port);
   mult_125_G2_FS_1_U1_0_4_0 : nand2 port map( a => n5826, b => n5827, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_4_0_port);
   mult_125_G2_FS_1_U5_0_3_3 : oai12 port map( b => n5824, c => n5825, a => 
                           mult_125_G2_FS_1_G_n_int_0_3_3_port, outb => 
                           mult_125_G2_FS_1_G_1_0_3_port);
   mult_125_G2_FS_1_U3_C_0_3_3 : xor2 port map( a => 
                           mult_125_G2_FS_1_PG_int_0_3_3_port, b => 
                           mult_125_G2_FS_1_C_1_3_3_port, outb => 
                           multiplier_sigs_1_17_port);
   mult_125_G2_FS_1_U3_B_0_3_3 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_3_3_port, b => 
                           mult_125_G2_FS_1_P_0_3_3_port, outb => n5823);
   mult_125_G2_FS_1_U2_0_3_3 : nand2 port map( a => mult_125_G2_A1_15_port, b 
                           => mult_125_G2_A2_15_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_3_3_port);
   mult_125_G2_FS_1_U1_0_3_3 : nand2 port map( a => n5821, b => n5822, outb => 
                           mult_125_G2_FS_1_P_0_3_3_port);
   mult_125_G2_FS_1_U3_B_0_3_2 : nand2 port map( a => 
                           mult_125_G2_FS_1_G_n_int_0_3_2_port, b => 
                           mult_125_G2_FS_1_P_0_3_2_port, outb => n5820);
   mult_125_G2_FS_1_U2_0_3_2 : nand2 port map( a => mult_125_G2_A1_14_port, b 
                           => mult_125_G2_A2_14_port, outb => 
                           mult_125_G2_FS_1_G_n_int_0_3_2_port);
   mult_125_G2_FS_1_U1_0_3_2 : nand2 port map( a => n5818, b => n5819, outb => 
                           mult_125_G2_FS_1_P_0_3_2_port);
   mult_125_G2_AN1_15 : inv port map( inb => coefficient_mem_array_1_15_port, 
                           outb => mult_125_G2_A_not_15_port);
   mult_125_G2_AN1_14 : inv port map( inb => coefficient_mem_array_1_14_port, 
                           outb => mult_125_G2_A_not_14_port);
   mult_125_G2_AN1_13 : inv port map( inb => coefficient_mem_array_1_13_port, 
                           outb => mult_125_G2_A_not_13_port);
   mult_125_G2_AN1_12 : inv port map( inb => coefficient_mem_array_1_12_port, 
                           outb => mult_125_G2_A_not_12_port);
   mult_125_G2_AN1_11 : inv port map( inb => coefficient_mem_array_1_11_port, 
                           outb => mult_125_G2_A_not_11_port);
   mult_125_G2_AN1_10 : inv port map( inb => coefficient_mem_array_1_10_port, 
                           outb => mult_125_G2_A_not_10_port);
   mult_125_G2_AN1_9 : inv port map( inb => coefficient_mem_array_1_9_port, 
                           outb => mult_125_G2_A_not_9_port);
   mult_125_G2_AN1_8 : inv port map( inb => coefficient_mem_array_1_8_port, 
                           outb => mult_125_G2_A_not_8_port);
   mult_125_G2_AN1_7 : inv port map( inb => coefficient_mem_array_1_7_port, 
                           outb => mult_125_G2_A_not_7_port);
   mult_125_G2_AN1_6 : inv port map( inb => coefficient_mem_array_1_6_port, 
                           outb => mult_125_G2_A_not_6_port);
   mult_125_G2_AN1_5 : inv port map( inb => coefficient_mem_array_1_5_port, 
                           outb => mult_125_G2_A_not_5_port);
   mult_125_G2_AN1_4 : inv port map( inb => coefficient_mem_array_1_4_port, 
                           outb => mult_125_G2_A_not_4_port);
   mult_125_G2_AN1_3 : inv port map( inb => coefficient_mem_array_1_3_port, 
                           outb => mult_125_G2_A_not_3_port);
   mult_125_G2_AN1_2 : inv port map( inb => coefficient_mem_array_1_2_port, 
                           outb => mult_125_G2_A_not_2_port);
   mult_125_G2_AN1_1 : inv port map( inb => coefficient_mem_array_1_1_port, 
                           outb => mult_125_G2_A_not_1_port);
   mult_125_G2_AN1_0 : inv port map( inb => coefficient_mem_array_1_0_port, 
                           outb => mult_125_G2_A_not_0_port);
   mult_125_G2_AN1_15_0 : inv port map( inb => input_sample_mem_15_port, outb 
                           => mult_125_G2_B_not_15_port);
   mult_125_G2_AN1_14_0 : inv port map( inb => input_sample_mem_14_port, outb 
                           => mult_125_G2_B_not_14_port);
   mult_125_G2_AN1_13_0 : inv port map( inb => input_sample_mem_13_port, outb 
                           => mult_125_G2_B_not_13_port);
   mult_125_G2_AN1_12_0 : inv port map( inb => input_sample_mem_12_port, outb 
                           => mult_125_G2_B_not_12_port);
   mult_125_G2_AN1_11_0 : inv port map( inb => input_sample_mem_11_port, outb 
                           => mult_125_G2_B_not_11_port);
   mult_125_G2_AN1_10_0 : inv port map( inb => input_sample_mem_10_port, outb 
                           => mult_125_G2_B_not_10_port);
   mult_125_G2_AN1_9_0 : inv port map( inb => input_sample_mem_9_port, outb => 
                           mult_125_G2_B_not_9_port);
   mult_125_G2_AN1_8_0 : inv port map( inb => input_sample_mem_8_port, outb => 
                           mult_125_G2_B_not_8_port);
   mult_125_G2_AN1_7_0 : inv port map( inb => input_sample_mem_7_port, outb => 
                           mult_125_G2_B_not_7_port);
   mult_125_G2_AN1_6_0 : inv port map( inb => input_sample_mem_6_port, outb => 
                           mult_125_G2_B_not_6_port);
   mult_125_G2_AN1_5_0 : inv port map( inb => input_sample_mem_5_port, outb => 
                           mult_125_G2_B_not_5_port);
   mult_125_G2_AN1_4_0 : inv port map( inb => input_sample_mem_4_port, outb => 
                           mult_125_G2_B_not_4_port);
   mult_125_G2_AN1_3_0 : inv port map( inb => input_sample_mem_3_port, outb => 
                           mult_125_G2_B_not_3_port);
   mult_125_G2_AN1_2_0 : inv port map( inb => input_sample_mem_2_port, outb => 
                           mult_125_G2_B_not_2_port);
   mult_125_G2_AN1_1_0 : inv port map( inb => input_sample_mem_1_port, outb => 
                           mult_125_G2_B_not_1_port);
   mult_125_G2_AN1_0_0 : inv port map( inb => input_sample_mem_0_port, outb => 
                           mult_125_G2_B_not_0_port);
   mult_125_G2_AN1_15_15 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_15_15_port);
   mult_125_G2_AN3_15_14 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_14_port, outb => 
                           mult_125_G2_ab_15_14_port);
   mult_125_G2_AN3_15_13 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_13_port, outb => 
                           mult_125_G2_ab_15_13_port);
   mult_125_G2_AN3_15_12 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_12_port, outb => 
                           mult_125_G2_ab_15_12_port);
   mult_125_G2_AN3_15_11 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_11_port, outb => 
                           mult_125_G2_ab_15_11_port);
   mult_125_G2_AN3_15_10 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_10_port, outb => 
                           mult_125_G2_ab_15_10_port);
   mult_125_G2_AN3_15_9 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_9_port, outb => 
                           mult_125_G2_ab_15_9_port);
   mult_125_G2_AN3_15_8 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_8_port, outb => 
                           mult_125_G2_ab_15_8_port);
   mult_125_G2_AN3_15_7 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_7_port, outb => 
                           mult_125_G2_ab_15_7_port);
   mult_125_G2_AN3_15_6 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_6_port, outb => 
                           mult_125_G2_ab_15_6_port);
   mult_125_G2_AN3_15_5 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_5_port, outb => 
                           mult_125_G2_ab_15_5_port);
   mult_125_G2_AN3_15_4 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_4_port, outb => 
                           mult_125_G2_ab_15_4_port);
   mult_125_G2_AN3_15_3 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_3_port, outb => 
                           mult_125_G2_ab_15_3_port);
   mult_125_G2_AN3_15_2 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_2_port, outb => 
                           mult_125_G2_ab_15_2_port);
   mult_125_G2_AN3_15_1 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_1_port, outb => 
                           mult_125_G2_ab_15_1_port);
   mult_125_G2_AN3_15_0 : nor2 port map( a => mult_125_G2_A_not_15_port, b => 
                           mult_125_G2_B_notx_0_port, outb => 
                           mult_125_G2_ab_15_0_port);
   mult_125_G2_AN2_14_15 : nor2 port map( a => mult_125_G2_A_notx_14_port, b =>
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_14_15_port);
   mult_125_G2_AN1_14_14 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_14_14_port);
   mult_125_G2_AN1_14_13 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_14_13_port);
   mult_125_G2_AN1_14_12 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_14_12_port);
   mult_125_G2_AN1_14_11 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_14_11_port);
   mult_125_G2_AN1_14_10 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_14_10_port);
   mult_125_G2_AN1_14_9 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_14_9_port);
   mult_125_G2_AN1_14_8 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_14_8_port);
   mult_125_G2_AN1_14_7 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_14_7_port);
   mult_125_G2_AN1_14_6 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_14_6_port);
   mult_125_G2_AN1_14_5 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_14_5_port);
   mult_125_G2_AN1_14_4 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_14_4_port);
   mult_125_G2_AN1_14_3 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_14_3_port);
   mult_125_G2_AN1_14_2 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_14_2_port);
   mult_125_G2_AN1_14_1 : nor2 port map( a => mult_125_G2_A_not_14_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_14_1_port);
   mult_125_G2_AN1_14_0_0 : nor2 port map( a => mult_125_G2_A_not_14_port, b =>
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_14_0_port);
   mult_125_G2_AN2_13_15 : nor2 port map( a => mult_125_G2_A_notx_13_port, b =>
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_13_15_port);
   mult_125_G2_AN1_13_14 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_13_14_port);
   mult_125_G2_AN1_13_13 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_13_13_port);
   mult_125_G2_AN1_13_12 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_13_12_port);
   mult_125_G2_AN1_13_11 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_13_11_port);
   mult_125_G2_AN1_13_10 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_13_10_port);
   mult_125_G2_AN1_13_9 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_13_9_port);
   mult_125_G2_AN1_13_8 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_13_8_port);
   mult_125_G2_AN1_13_7 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_13_7_port);
   mult_125_G2_AN1_13_6 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_13_6_port);
   mult_125_G2_AN1_13_5 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_13_5_port);
   mult_125_G2_AN1_13_4 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_13_4_port);
   mult_125_G2_AN1_13_3 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_13_3_port);
   mult_125_G2_AN1_13_2 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_13_2_port);
   mult_125_G2_AN1_13_1 : nor2 port map( a => mult_125_G2_A_not_13_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_13_1_port);
   mult_125_G2_AN1_13_0_0 : nor2 port map( a => mult_125_G2_A_not_13_port, b =>
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_13_0_port);
   mult_125_G2_AN2_12_15 : nor2 port map( a => mult_125_G2_A_notx_12_port, b =>
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_12_15_port);
   mult_125_G2_AN1_12_14 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_12_14_port);
   mult_125_G2_AN1_12_13 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_12_13_port);
   mult_125_G2_AN1_12_12 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_12_12_port);
   mult_125_G2_AN1_12_11 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_12_11_port);
   mult_125_G2_AN1_12_10 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_12_10_port);
   mult_125_G2_AN1_12_9 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_12_9_port);
   mult_125_G2_AN1_12_8 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_12_8_port);
   mult_125_G2_AN1_12_7 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_12_7_port);
   mult_125_G2_AN1_12_6 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_12_6_port);
   mult_125_G2_AN1_12_5 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_12_5_port);
   mult_125_G2_AN1_12_4 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_12_4_port);
   mult_125_G2_AN1_12_3 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_12_3_port);
   mult_125_G2_AN1_12_2 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_12_2_port);
   mult_125_G2_AN1_12_1 : nor2 port map( a => mult_125_G2_A_not_12_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_12_1_port);
   mult_125_G2_AN1_12_0_0 : nor2 port map( a => mult_125_G2_A_not_12_port, b =>
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_12_0_port);
   mult_125_G2_AN2_11_15 : nor2 port map( a => mult_125_G2_A_notx_11_port, b =>
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_11_15_port);
   mult_125_G2_AN1_11_14 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_11_14_port);
   mult_125_G2_AN1_11_13 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_11_13_port);
   mult_125_G2_AN1_11_12 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_11_12_port);
   mult_125_G2_AN1_11_11 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_11_11_port);
   mult_125_G2_AN1_11_10 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_11_10_port);
   mult_125_G2_AN1_11_9 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_11_9_port);
   mult_125_G2_AN1_11_8 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_11_8_port);
   mult_125_G2_AN1_11_7 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_11_7_port);
   mult_125_G2_AN1_11_6 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_11_6_port);
   mult_125_G2_AN1_11_5 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_11_5_port);
   mult_125_G2_AN1_11_4 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_11_4_port);
   mult_125_G2_AN1_11_3 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_11_3_port);
   mult_125_G2_AN1_11_2 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_11_2_port);
   mult_125_G2_AN1_11_1 : nor2 port map( a => mult_125_G2_A_not_11_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_11_1_port);
   mult_125_G2_AN1_11_0_0 : nor2 port map( a => mult_125_G2_A_not_11_port, b =>
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_11_0_port);
   mult_125_G2_AN2_10_15 : nor2 port map( a => mult_125_G2_A_notx_10_port, b =>
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_10_15_port);
   mult_125_G2_AN1_10_14 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_10_14_port);
   mult_125_G2_AN1_10_13 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_10_13_port);
   mult_125_G2_AN1_10_12 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_10_12_port);
   mult_125_G2_AN1_10_11 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_10_11_port);
   mult_125_G2_AN1_10_10 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_10_10_port);
   mult_125_G2_AN1_10_9 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_10_9_port);
   mult_125_G2_AN1_10_8 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_10_8_port);
   mult_125_G2_AN1_10_7 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_10_7_port);
   mult_125_G2_AN1_10_6 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_10_6_port);
   mult_125_G2_AN1_10_5 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_10_5_port);
   mult_125_G2_AN1_10_4 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_10_4_port);
   mult_125_G2_AN1_10_3 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_10_3_port);
   mult_125_G2_AN1_10_2 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_10_2_port);
   mult_125_G2_AN1_10_1 : nor2 port map( a => mult_125_G2_A_not_10_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_10_1_port);
   mult_125_G2_AN1_10_0_0 : nor2 port map( a => mult_125_G2_A_not_10_port, b =>
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_10_0_port);
   mult_125_G2_AN2_9_15 : nor2 port map( a => mult_125_G2_A_notx_9_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_9_15_port);
   mult_125_G2_AN1_9_14 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_9_14_port);
   mult_125_G2_AN1_9_13 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_9_13_port);
   mult_125_G2_AN1_9_12 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_9_12_port);
   mult_125_G2_AN1_9_11 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_9_11_port);
   mult_125_G2_AN1_9_10 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_9_10_port);
   mult_125_G2_AN1_9_9 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_9_9_port);
   mult_125_G2_AN1_9_8 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_9_8_port);
   mult_125_G2_AN1_9_7 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_9_7_port);
   mult_125_G2_AN1_9_6 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_9_6_port);
   mult_125_G2_AN1_9_5 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_9_5_port);
   mult_125_G2_AN1_9_4 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_9_4_port);
   mult_125_G2_AN1_9_3 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_9_3_port);
   mult_125_G2_AN1_9_2 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_9_2_port);
   mult_125_G2_AN1_9_1 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_9_1_port);
   mult_125_G2_AN1_9_0_0 : nor2 port map( a => mult_125_G2_A_not_9_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_9_0_port);
   mult_125_G2_AN2_8_15 : nor2 port map( a => mult_125_G2_A_notx_8_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_8_15_port);
   mult_125_G2_AN1_8_14 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_8_14_port);
   mult_125_G2_AN1_8_13 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_8_13_port);
   mult_125_G2_AN1_8_12 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_8_12_port);
   mult_125_G2_AN1_8_11 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_8_11_port);
   mult_125_G2_AN1_8_10 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_8_10_port);
   mult_125_G2_AN1_8_9 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_8_9_port);
   mult_125_G2_AN1_8_8 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_8_8_port);
   mult_125_G2_AN1_8_7 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_8_7_port);
   mult_125_G2_AN1_8_6 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_8_6_port);
   mult_125_G2_AN1_8_5 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_8_5_port);
   mult_125_G2_AN1_8_4 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_8_4_port);
   mult_125_G2_AN1_8_3 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_8_3_port);
   mult_125_G2_AN1_8_2 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_8_2_port);
   mult_125_G2_AN1_8_1 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_8_1_port);
   mult_125_G2_AN1_8_0_0 : nor2 port map( a => mult_125_G2_A_not_8_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_8_0_port);
   mult_125_G2_AN2_7_15 : nor2 port map( a => mult_125_G2_A_notx_7_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_7_15_port);
   mult_125_G2_AN1_7_14 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_7_14_port);
   mult_125_G2_AN1_7_13 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_7_13_port);
   mult_125_G2_AN1_7_12 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_7_12_port);
   mult_125_G2_AN1_7_11 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_7_11_port);
   mult_125_G2_AN1_7_10 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_7_10_port);
   mult_125_G2_AN1_7_9 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_7_9_port);
   mult_125_G2_AN1_7_8 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_7_8_port);
   mult_125_G2_AN1_7_7 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_7_7_port);
   mult_125_G2_AN1_7_6 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_7_6_port);
   mult_125_G2_AN1_7_5 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_7_5_port);
   mult_125_G2_AN1_7_4 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_7_4_port);
   mult_125_G2_AN1_7_3 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_7_3_port);
   mult_125_G2_AN1_7_2 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_7_2_port);
   mult_125_G2_AN1_7_1 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_7_1_port);
   mult_125_G2_AN1_7_0_0 : nor2 port map( a => mult_125_G2_A_not_7_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_7_0_port);
   mult_125_G2_AN2_6_15 : nor2 port map( a => mult_125_G2_A_notx_6_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_6_15_port);
   mult_125_G2_AN1_6_14 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_6_14_port);
   mult_125_G2_AN1_6_13 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_6_13_port);
   mult_125_G2_AN1_6_12 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_6_12_port);
   mult_125_G2_AN1_6_11 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_6_11_port);
   mult_125_G2_AN1_6_10 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_6_10_port);
   mult_125_G2_AN1_6_9 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_6_9_port);
   mult_125_G2_AN1_6_8 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_6_8_port);
   mult_125_G2_AN1_6_7 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_6_7_port);
   mult_125_G2_AN1_6_6 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_6_6_port);
   mult_125_G2_AN1_6_5 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_6_5_port);
   mult_125_G2_AN1_6_4 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_6_4_port);
   mult_125_G2_AN1_6_3 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_6_3_port);
   mult_125_G2_AN1_6_2 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_6_2_port);
   mult_125_G2_AN1_6_1 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_6_1_port);
   mult_125_G2_AN1_6_0_0 : nor2 port map( a => mult_125_G2_A_not_6_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_6_0_port);
   mult_125_G2_AN2_5_15 : nor2 port map( a => mult_125_G2_A_notx_5_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_5_15_port);
   mult_125_G2_AN1_5_14 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_5_14_port);
   mult_125_G2_AN1_5_13 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_5_13_port);
   mult_125_G2_AN1_5_12 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_5_12_port);
   mult_125_G2_AN1_5_11 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_5_11_port);
   mult_125_G2_AN1_5_10 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_5_10_port);
   mult_125_G2_AN1_5_9 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_5_9_port);
   mult_125_G2_AN1_5_8 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_5_8_port);
   mult_125_G2_AN1_5_7 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_5_7_port);
   mult_125_G2_AN1_5_6 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_5_6_port);
   mult_125_G2_AN1_5_5 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_5_5_port);
   mult_125_G2_AN1_5_4 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_5_4_port);
   mult_125_G2_AN1_5_3 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_5_3_port);
   mult_125_G2_AN1_5_2 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_5_2_port);
   mult_125_G2_AN1_5_1 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_5_1_port);
   mult_125_G2_AN1_5_0_0 : nor2 port map( a => mult_125_G2_A_not_5_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_5_0_port);
   mult_125_G2_AN2_4_15 : nor2 port map( a => mult_125_G2_A_notx_4_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_4_15_port);
   mult_125_G2_AN1_4_14 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_4_14_port);
   mult_125_G2_AN1_4_13 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_4_13_port);
   mult_125_G2_AN1_4_12 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_4_12_port);
   mult_125_G2_AN1_4_11 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_4_11_port);
   mult_125_G2_AN1_4_10 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_4_10_port);
   mult_125_G2_AN1_4_9 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_4_9_port);
   mult_125_G2_AN1_4_8 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_4_8_port);
   mult_125_G2_AN1_4_7 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_4_7_port);
   mult_125_G2_AN1_4_6 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_4_6_port);
   mult_125_G2_AN1_4_5 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_4_5_port);
   mult_125_G2_AN1_4_4 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_4_4_port);
   mult_125_G2_AN1_4_3 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_4_3_port);
   mult_125_G2_AN1_4_2 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_4_2_port);
   mult_125_G2_AN1_4_1 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_4_1_port);
   mult_125_G2_AN1_4_0_0 : nor2 port map( a => mult_125_G2_A_not_4_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_4_0_port);
   mult_125_G2_AN2_3_15 : nor2 port map( a => mult_125_G2_A_notx_3_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_3_15_port);
   mult_125_G2_AN1_3_14 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_3_14_port);
   mult_125_G2_AN1_3_13 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_3_13_port);
   mult_125_G2_AN1_3_12 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_3_12_port);
   mult_125_G2_AN1_3_11 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_3_11_port);
   mult_125_G2_AN1_3_10 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_3_10_port);
   mult_125_G2_AN1_3_9 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_3_9_port);
   mult_125_G2_AN1_3_8 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_3_8_port);
   mult_125_G2_AN1_3_7 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_3_7_port);
   mult_125_G2_AN1_3_6 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_3_6_port);
   mult_125_G2_AN1_3_5 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_3_5_port);
   mult_125_G2_AN1_3_4 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_3_4_port);
   mult_125_G2_AN1_3_3 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_3_3_port);
   mult_125_G2_AN1_3_2 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_3_2_port);
   mult_125_G2_AN1_3_1 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_3_1_port);
   mult_125_G2_AN1_3_0_0 : nor2 port map( a => mult_125_G2_A_not_3_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_3_0_port);
   mult_125_G2_AN2_2_15 : nor2 port map( a => mult_125_G2_A_notx_2_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_2_15_port);
   mult_125_G2_AN1_2_14 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_2_14_port);
   mult_125_G2_AN1_2_13 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_2_13_port);
   mult_125_G2_AN1_2_12 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_2_12_port);
   mult_125_G2_AN1_2_11 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_2_11_port);
   mult_125_G2_AN1_2_10 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_2_10_port);
   mult_125_G2_AN1_2_9 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_2_9_port);
   mult_125_G2_AN1_2_8 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_2_8_port);
   mult_125_G2_AN1_2_7 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_2_7_port);
   mult_125_G2_AN1_2_6 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_2_6_port);
   mult_125_G2_AN1_2_5 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_2_5_port);
   mult_125_G2_AN1_2_4 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_2_4_port);
   mult_125_G2_AN1_2_3 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_2_3_port);
   mult_125_G2_AN1_2_2 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_2_2_port);
   mult_125_G2_AN1_2_1 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_2_1_port);
   mult_125_G2_AN1_2_0_0 : nor2 port map( a => mult_125_G2_A_not_2_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_2_0_port);
   mult_125_G2_AN2_1_15 : nor2 port map( a => mult_125_G2_A_notx_1_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_1_15_port);
   mult_125_G2_AN1_1_14 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_1_14_port);
   mult_125_G2_AN1_1_13 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_1_13_port);
   mult_125_G2_AN1_1_12 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_1_12_port);
   mult_125_G2_AN1_1_11 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_1_11_port);
   mult_125_G2_AN1_1_10 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_1_10_port);
   mult_125_G2_AN1_1_9 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_1_9_port);
   mult_125_G2_AN1_1_8 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_1_8_port);
   mult_125_G2_AN1_1_7 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_1_7_port);
   mult_125_G2_AN1_1_6 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_1_6_port);
   mult_125_G2_AN1_1_5 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_1_5_port);
   mult_125_G2_AN1_1_4 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_1_4_port);
   mult_125_G2_AN1_1_3 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_1_3_port);
   mult_125_G2_AN1_1_2 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_1_2_port);
   mult_125_G2_AN1_1_1 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_1_1_port);
   mult_125_G2_AN1_1_0_0 : nor2 port map( a => mult_125_G2_A_not_1_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_ab_1_0_port);
   mult_125_G2_AN2_0_15 : nor2 port map( a => mult_125_G2_A_notx_0_port, b => 
                           mult_125_G2_B_not_15_port, outb => 
                           mult_125_G2_ab_0_15_port);
   mult_125_G2_AN1_0_14 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_ab_0_14_port);
   mult_125_G2_AN1_0_13 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_ab_0_13_port);
   mult_125_G2_AN1_0_12 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_ab_0_12_port);
   mult_125_G2_AN1_0_11 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_ab_0_11_port);
   mult_125_G2_AN1_0_10 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_ab_0_10_port);
   mult_125_G2_AN1_0_9 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_ab_0_9_port);
   mult_125_G2_AN1_0_8 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_ab_0_8_port);
   mult_125_G2_AN1_0_7 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_ab_0_7_port);
   mult_125_G2_AN1_0_6 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_ab_0_6_port);
   mult_125_G2_AN1_0_5 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_ab_0_5_port);
   mult_125_G2_AN1_0_4 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_ab_0_4_port);
   mult_125_G2_AN1_0_3 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_ab_0_3_port);
   mult_125_G2_AN1_0_2 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_ab_0_2_port);
   mult_125_G2_AN1_0_1 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_ab_0_1_port);
   mult_125_G2_AN1_0_0_0 : nor2 port map( a => mult_125_G2_A_not_0_port, b => 
                           mult_125_G2_B_not_0_port, outb => 
                           multiplier_sigs_1_0_port);
   mult_125_FS_1_U6_1_1_3 : oai12 port map( b => n5782, c => n5783, a => n5784,
                           outb => mult_125_FS_1_C_1_7_0_port);
   mult_125_FS_1_U6_1_1_2 : oai12 port map( b => n5779, c => n5780, a => n5781,
                           outb => mult_125_FS_1_C_1_6_0_port);
   mult_125_FS_1_U6_1_1_1 : oai12 port map( b => n5776, c => n5777, a => n5778,
                           outb => mult_125_FS_1_C_1_5_0_port);
   mult_125_FS_1_U6_0_7_1 : oai12 port map( b => n5773, c => n5774, a => 
                           mult_125_FS_1_G_n_int_0_7_0_port, outb => 
                           mult_125_FS_1_C_1_7_1_port);
   mult_125_FS_1_U3_C_0_7_1 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_7_1_port, b => 
                           mult_125_FS_1_C_1_7_1_port, outb => 
                           multiplier_sigs_0_31_port);
   mult_125_FS_1_U3_B_0_7_1 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_7_1_port, b => 
                           mult_125_FS_1_P_0_7_1_port, outb => n5772);
   mult_125_FS_1_U2_0_7_1 : nand2 port map( a => mult_125_A1_29_port, b => 
                           mult_125_A2_29_port, outb => 
                           mult_125_FS_1_G_n_int_0_7_1_port);
   mult_125_FS_1_U1_0_7_1 : nand2 port map( a => n5770, b => n5771, outb => 
                           mult_125_FS_1_P_0_7_1_port);
   mult_125_FS_1_U3_C_0_7_0 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_7_0_port, b => 
                           mult_125_FS_1_C_1_7_0_port, outb => 
                           multiplier_sigs_0_30_port);
   mult_125_FS_1_U3_B_0_7_0 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_7_0_port, b => 
                           mult_125_FS_1_TEMP_P_0_7_0_port, outb => n5769);
   mult_125_FS_1_U2_0_7_0 : nand2 port map( a => mult_125_A1_28_port, b => 
                           mult_125_A2_28_port, outb => 
                           mult_125_FS_1_G_n_int_0_7_0_port);
   mult_125_FS_1_U1_0_7_0 : nand2 port map( a => n5767, b => n5768, outb => 
                           mult_125_FS_1_TEMP_P_0_7_0_port);
   mult_125_FS_1_U6_0_6_3 : oai12 port map( b => n5765, c => n5766, a => 
                           mult_125_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_FS_1_C_1_6_3_port);
   mult_125_FS_1_U5_0_6_3 : oai12 port map( b => n5763, c => n5764, a => 
                           mult_125_FS_1_G_n_int_0_6_3_port, outb => 
                           mult_125_FS_1_G_1_1_2_port);
   mult_125_FS_1_U4_0_6_3 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_6_2_port, b => 
                           mult_125_FS_1_P_0_6_3_port, outb => n5783);
   mult_125_FS_1_U3_C_0_6_3 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_6_3_port, b => 
                           mult_125_FS_1_C_1_6_3_port, outb => 
                           multiplier_sigs_0_29_port);
   mult_125_FS_1_U3_B_0_6_3 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_6_3_port, b => 
                           mult_125_FS_1_P_0_6_3_port, outb => n5762);
   mult_125_FS_1_U2_0_6_3 : nand2 port map( a => mult_125_A1_27_port, b => 
                           mult_125_A2_27_port, outb => 
                           mult_125_FS_1_G_n_int_0_6_3_port);
   mult_125_FS_1_U1_0_6_3 : nand2 port map( a => n5760, b => n5761, outb => 
                           mult_125_FS_1_P_0_6_3_port);
   mult_125_FS_1_U6_0_6_2 : oai12 port map( b => n5758, c => n5759, a => 
                           mult_125_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_FS_1_C_1_6_2_port);
   mult_125_FS_1_U5_0_6_2 : oai12 port map( b => n5757, c => n5766, a => 
                           mult_125_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_FS_1_TEMP_G_0_6_2_port);
   mult_125_FS_1_U4_0_6_2 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_6_1_port, b => 
                           mult_125_FS_1_P_0_6_2_port, outb => n5756);
   mult_125_FS_1_U3_C_0_6_2 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_6_2_port, b => 
                           mult_125_FS_1_C_1_6_2_port, outb => 
                           multiplier_sigs_0_28_port);
   mult_125_FS_1_U3_B_0_6_2 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_6_2_port, b => 
                           mult_125_FS_1_P_0_6_2_port, outb => n5755);
   mult_125_FS_1_U2_0_6_2 : nand2 port map( a => mult_125_A1_26_port, b => 
                           mult_125_A2_26_port, outb => 
                           mult_125_FS_1_G_n_int_0_6_2_port);
   mult_125_FS_1_U1_0_6_2 : nand2 port map( a => n5753, b => n5754, outb => 
                           mult_125_FS_1_P_0_6_2_port);
   mult_125_FS_1_U6_0_6_1 : oai12 port map( b => n5782, c => n5752, a => 
                           mult_125_FS_1_G_n_int_0_6_0_port, outb => 
                           mult_125_FS_1_C_1_6_1_port);
   mult_125_FS_1_U5_0_6_1 : oai12 port map( b => 
                           mult_125_FS_1_G_n_int_0_6_0_port, c => n5759, a => 
                           mult_125_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_FS_1_TEMP_G_0_6_1_port);
   mult_125_FS_1_U4_0_6_1 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_6_0_port, b => 
                           mult_125_FS_1_P_0_6_1_port, outb => n5751);
   mult_125_FS_1_U3_C_0_6_1 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_6_1_port, b => 
                           mult_125_FS_1_C_1_6_1_port, outb => 
                           multiplier_sigs_0_27_port);
   mult_125_FS_1_U3_B_0_6_1 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_6_1_port, b => 
                           mult_125_FS_1_P_0_6_1_port, outb => n5750);
   mult_125_FS_1_U2_0_6_1 : nand2 port map( a => mult_125_A1_25_port, b => 
                           mult_125_A2_25_port, outb => 
                           mult_125_FS_1_G_n_int_0_6_1_port);
   mult_125_FS_1_U1_0_6_1 : nand2 port map( a => n5748, b => n5749, outb => 
                           mult_125_FS_1_P_0_6_1_port);
   mult_125_FS_1_U3_C_0_6_0 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_6_0_port, b => 
                           mult_125_FS_1_C_1_6_0_port, outb => 
                           multiplier_sigs_0_26_port);
   mult_125_FS_1_U3_B_0_6_0 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_6_0_port, b => 
                           mult_125_FS_1_TEMP_P_0_6_0_port, outb => n5747);
   mult_125_FS_1_U2_0_6_0 : nand2 port map( a => mult_125_A1_24_port, b => 
                           mult_125_A2_24_port, outb => 
                           mult_125_FS_1_G_n_int_0_6_0_port);
   mult_125_FS_1_U1_0_6_0 : nand2 port map( a => n5745, b => n5746, outb => 
                           mult_125_FS_1_TEMP_P_0_6_0_port);
   mult_125_FS_1_U6_0_5_3 : oai12 port map( b => n5743, c => n5744, a => 
                           mult_125_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_FS_1_C_1_5_3_port);
   mult_125_FS_1_U5_0_5_3 : oai12 port map( b => n5741, c => n5742, a => 
                           mult_125_FS_1_G_n_int_0_5_3_port, outb => 
                           mult_125_FS_1_G_1_1_1_port);
   mult_125_FS_1_U4_0_5_3 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_5_2_port, b => 
                           mult_125_FS_1_P_0_5_3_port, outb => n5780);
   mult_125_FS_1_U3_C_0_5_3 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_5_3_port, b => 
                           mult_125_FS_1_C_1_5_3_port, outb => 
                           multiplier_sigs_0_25_port);
   mult_125_FS_1_U3_B_0_5_3 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_5_3_port, b => 
                           mult_125_FS_1_P_0_5_3_port, outb => n5740);
   mult_125_FS_1_U2_0_5_3 : nand2 port map( a => mult_125_A1_23_port, b => 
                           mult_125_A2_23_port, outb => 
                           mult_125_FS_1_G_n_int_0_5_3_port);
   mult_125_FS_1_U1_0_5_3 : nand2 port map( a => n5738, b => n5739, outb => 
                           mult_125_FS_1_P_0_5_3_port);
   mult_125_FS_1_U6_0_5_2 : oai12 port map( b => n5736, c => n5737, a => 
                           mult_125_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_FS_1_C_1_5_2_port);
   mult_125_FS_1_U5_0_5_2 : oai12 port map( b => n5735, c => n5744, a => 
                           mult_125_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_FS_1_TEMP_G_0_5_2_port);
   mult_125_FS_1_U4_0_5_2 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_5_1_port, b => 
                           mult_125_FS_1_P_0_5_2_port, outb => n5734);
   mult_125_FS_1_U3_C_0_5_2 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_5_2_port, b => 
                           mult_125_FS_1_C_1_5_2_port, outb => 
                           multiplier_sigs_0_24_port);
   mult_125_FS_1_U3_B_0_5_2 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_5_2_port, b => 
                           mult_125_FS_1_P_0_5_2_port, outb => n5733);
   mult_125_FS_1_U2_0_5_2 : nand2 port map( a => mult_125_A1_22_port, b => 
                           mult_125_A2_22_port, outb => 
                           mult_125_FS_1_G_n_int_0_5_2_port);
   mult_125_FS_1_U1_0_5_2 : nand2 port map( a => n5731, b => n5732, outb => 
                           mult_125_FS_1_P_0_5_2_port);
   mult_125_FS_1_U6_0_5_1 : oai12 port map( b => n5779, c => n5730, a => 
                           mult_125_FS_1_G_n_int_0_5_0_port, outb => 
                           mult_125_FS_1_C_1_5_1_port);
   mult_125_FS_1_U5_0_5_1 : oai12 port map( b => 
                           mult_125_FS_1_G_n_int_0_5_0_port, c => n5737, a => 
                           mult_125_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_FS_1_TEMP_G_0_5_1_port);
   mult_125_FS_1_U4_0_5_1 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_5_0_port, b => 
                           mult_125_FS_1_P_0_5_1_port, outb => n5729);
   mult_125_FS_1_U3_C_0_5_1 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_5_1_port, b => 
                           mult_125_FS_1_C_1_5_1_port, outb => 
                           multiplier_sigs_0_23_port);
   mult_125_FS_1_U3_B_0_5_1 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_5_1_port, b => 
                           mult_125_FS_1_P_0_5_1_port, outb => n5728);
   mult_125_FS_1_U2_0_5_1 : nand2 port map( a => mult_125_A1_21_port, b => 
                           mult_125_A2_21_port, outb => 
                           mult_125_FS_1_G_n_int_0_5_1_port);
   mult_125_FS_1_U1_0_5_1 : nand2 port map( a => n5726, b => n5727, outb => 
                           mult_125_FS_1_P_0_5_1_port);
   mult_125_FS_1_U3_C_0_5_0 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_5_0_port, b => 
                           mult_125_FS_1_C_1_5_0_port, outb => 
                           multiplier_sigs_0_22_port);
   mult_125_FS_1_U3_B_0_5_0 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_5_0_port, b => 
                           mult_125_FS_1_TEMP_P_0_5_0_port, outb => n5725);
   mult_125_FS_1_U2_0_5_0 : nand2 port map( a => mult_125_A1_20_port, b => 
                           mult_125_A2_20_port, outb => 
                           mult_125_FS_1_G_n_int_0_5_0_port);
   mult_125_FS_1_U1_0_5_0 : nand2 port map( a => n5723, b => n5724, outb => 
                           mult_125_FS_1_TEMP_P_0_5_0_port);
   mult_125_FS_1_U6_0_4_3 : oai12 port map( b => n5721, c => n5722, a => 
                           mult_125_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_FS_1_C_1_4_3_port);
   mult_125_FS_1_U5_0_4_3 : oai12 port map( b => n5719, c => n5720, a => 
                           mult_125_FS_1_G_n_int_0_4_3_port, outb => 
                           mult_125_FS_1_G_1_1_0_port);
   mult_125_FS_1_U4_0_4_3 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_4_2_port, b => 
                           mult_125_FS_1_P_0_4_3_port, outb => n5777);
   mult_125_FS_1_U3_C_0_4_3 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_4_3_port, b => 
                           mult_125_FS_1_C_1_4_3_port, outb => 
                           multiplier_sigs_0_21_port);
   mult_125_FS_1_U3_B_0_4_3 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_4_3_port, b => 
                           mult_125_FS_1_P_0_4_3_port, outb => n5718);
   mult_125_FS_1_U2_0_4_3 : nand2 port map( a => mult_125_A1_19_port, b => 
                           mult_125_A2_19_port, outb => 
                           mult_125_FS_1_G_n_int_0_4_3_port);
   mult_125_FS_1_U1_0_4_3 : nand2 port map( a => n5716, b => n5717, outb => 
                           mult_125_FS_1_P_0_4_3_port);
   mult_125_FS_1_U6_0_4_2 : oai12 port map( b => n5714, c => n5715, a => 
                           mult_125_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_FS_1_C_1_4_2_port);
   mult_125_FS_1_U5_0_4_2 : oai12 port map( b => n5713, c => n5722, a => 
                           mult_125_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_FS_1_TEMP_G_0_4_2_port);
   mult_125_FS_1_U4_0_4_2 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_4_1_port, b => 
                           mult_125_FS_1_P_0_4_2_port, outb => n5712);
   mult_125_FS_1_U3_C_0_4_2 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_4_2_port, b => 
                           mult_125_FS_1_C_1_4_2_port, outb => 
                           multiplier_sigs_0_20_port);
   mult_125_FS_1_U3_B_0_4_2 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_4_2_port, b => 
                           mult_125_FS_1_P_0_4_2_port, outb => n5711);
   mult_125_FS_1_U2_0_4_2 : nand2 port map( a => mult_125_A1_18_port, b => 
                           mult_125_A2_18_port, outb => 
                           mult_125_FS_1_G_n_int_0_4_2_port);
   mult_125_FS_1_U1_0_4_2 : nand2 port map( a => n5709, b => n5710, outb => 
                           mult_125_FS_1_P_0_4_2_port);
   mult_125_FS_1_U6_0_4_1 : oai12 port map( b => n5776, c => n5708, a => 
                           mult_125_FS_1_G_n_int_0_4_0_port, outb => 
                           mult_125_FS_1_C_1_4_1_port);
   mult_125_FS_1_U5_0_4_1 : oai12 port map( b => 
                           mult_125_FS_1_G_n_int_0_4_0_port, c => n5715, a => 
                           mult_125_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_FS_1_TEMP_G_0_4_1_port);
   mult_125_FS_1_U4_0_4_1 : nand2 port map( a => 
                           mult_125_FS_1_TEMP_P_0_4_0_port, b => 
                           mult_125_FS_1_P_0_4_1_port, outb => n5707);
   mult_125_FS_1_U3_C_0_4_1 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_4_1_port, b => 
                           mult_125_FS_1_C_1_4_1_port, outb => 
                           multiplier_sigs_0_19_port);
   mult_125_FS_1_U3_B_0_4_1 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_4_1_port, b => 
                           mult_125_FS_1_P_0_4_1_port, outb => n5706);
   mult_125_FS_1_U2_0_4_1 : nand2 port map( a => mult_125_A1_17_port, b => 
                           mult_125_A2_17_port, outb => 
                           mult_125_FS_1_G_n_int_0_4_1_port);
   mult_125_FS_1_U1_0_4_1 : nand2 port map( a => n5704, b => n5705, outb => 
                           mult_125_FS_1_P_0_4_1_port);
   mult_125_FS_1_U3_C_0_4_0 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_4_0_port, b => 
                           mult_125_FS_1_C_1_4_0_port, outb => 
                           multiplier_sigs_0_18_port);
   mult_125_FS_1_U3_B_0_4_0 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_4_0_port, b => 
                           mult_125_FS_1_TEMP_P_0_4_0_port, outb => n5703);
   mult_125_FS_1_U2_0_4_0 : nand2 port map( a => mult_125_A1_16_port, b => 
                           mult_125_A2_16_port, outb => 
                           mult_125_FS_1_G_n_int_0_4_0_port);
   mult_125_FS_1_U1_0_4_0 : nand2 port map( a => n5701, b => n5702, outb => 
                           mult_125_FS_1_TEMP_P_0_4_0_port);
   mult_125_FS_1_U5_0_3_3 : oai12 port map( b => n5699, c => n5700, a => 
                           mult_125_FS_1_G_n_int_0_3_3_port, outb => 
                           mult_125_FS_1_G_1_0_3_port);
   mult_125_FS_1_U3_C_0_3_3 : xor2 port map( a => 
                           mult_125_FS_1_PG_int_0_3_3_port, b => 
                           mult_125_FS_1_C_1_3_3_port, outb => 
                           multiplier_sigs_0_17_port);
   mult_125_FS_1_U3_B_0_3_3 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_3_3_port, b => 
                           mult_125_FS_1_P_0_3_3_port, outb => n5698);
   mult_125_FS_1_U2_0_3_3 : nand2 port map( a => mult_125_A1_15_port, b => 
                           mult_125_A2_15_port, outb => 
                           mult_125_FS_1_G_n_int_0_3_3_port);
   mult_125_FS_1_U1_0_3_3 : nand2 port map( a => n5696, b => n5697, outb => 
                           mult_125_FS_1_P_0_3_3_port);
   mult_125_FS_1_U3_B_0_3_2 : nand2 port map( a => 
                           mult_125_FS_1_G_n_int_0_3_2_port, b => 
                           mult_125_FS_1_P_0_3_2_port, outb => n5695);
   mult_125_FS_1_U2_0_3_2 : nand2 port map( a => mult_125_A1_14_port, b => 
                           mult_125_A2_14_port, outb => 
                           mult_125_FS_1_G_n_int_0_3_2_port);
   mult_125_FS_1_U1_0_3_2 : nand2 port map( a => n5693, b => n5694, outb => 
                           mult_125_FS_1_P_0_3_2_port);
   mult_125_AN1_15 : inv port map( inb => coefficient_mem_array_0_15_port, outb
                           => mult_125_A_not_15_port);
   mult_125_AN1_14 : inv port map( inb => coefficient_mem_array_0_14_port, outb
                           => mult_125_A_not_14_port);
   mult_125_AN1_13 : inv port map( inb => coefficient_mem_array_0_13_port, outb
                           => mult_125_A_not_13_port);
   mult_125_AN1_12 : inv port map( inb => coefficient_mem_array_0_12_port, outb
                           => mult_125_A_not_12_port);
   mult_125_AN1_11 : inv port map( inb => coefficient_mem_array_0_11_port, outb
                           => mult_125_A_not_11_port);
   mult_125_AN1_10 : inv port map( inb => coefficient_mem_array_0_10_port, outb
                           => mult_125_A_not_10_port);
   mult_125_AN1_9 : inv port map( inb => coefficient_mem_array_0_9_port, outb 
                           => mult_125_A_not_9_port);
   mult_125_AN1_8 : inv port map( inb => coefficient_mem_array_0_8_port, outb 
                           => mult_125_A_not_8_port);
   mult_125_AN1_7 : inv port map( inb => coefficient_mem_array_0_7_port, outb 
                           => mult_125_A_not_7_port);
   mult_125_AN1_6 : inv port map( inb => coefficient_mem_array_0_6_port, outb 
                           => mult_125_A_not_6_port);
   mult_125_AN1_5 : inv port map( inb => coefficient_mem_array_0_5_port, outb 
                           => mult_125_A_not_5_port);
   mult_125_AN1_4 : inv port map( inb => coefficient_mem_array_0_4_port, outb 
                           => mult_125_A_not_4_port);
   mult_125_AN1_3 : inv port map( inb => coefficient_mem_array_0_3_port, outb 
                           => mult_125_A_not_3_port);
   mult_125_AN1_2 : inv port map( inb => coefficient_mem_array_0_2_port, outb 
                           => mult_125_A_not_2_port);
   mult_125_AN1_1 : inv port map( inb => coefficient_mem_array_0_1_port, outb 
                           => mult_125_A_not_1_port);
   mult_125_AN1_0 : inv port map( inb => coefficient_mem_array_0_0_port, outb 
                           => mult_125_A_not_0_port);
   mult_125_AN1_15_0 : inv port map( inb => input_sample_mem_15_port, outb => 
                           mult_125_B_not_15_port);
   mult_125_AN1_14_0 : inv port map( inb => input_sample_mem_14_port, outb => 
                           mult_125_B_not_14_port);
   mult_125_AN1_13_0 : inv port map( inb => input_sample_mem_13_port, outb => 
                           mult_125_B_not_13_port);
   mult_125_AN1_12_0 : inv port map( inb => input_sample_mem_12_port, outb => 
                           mult_125_B_not_12_port);
   mult_125_AN1_11_0 : inv port map( inb => input_sample_mem_11_port, outb => 
                           mult_125_B_not_11_port);
   mult_125_AN1_10_0 : inv port map( inb => input_sample_mem_10_port, outb => 
                           mult_125_B_not_10_port);
   mult_125_AN1_9_0 : inv port map( inb => input_sample_mem_9_port, outb => 
                           mult_125_B_not_9_port);
   mult_125_AN1_8_0 : inv port map( inb => input_sample_mem_8_port, outb => 
                           mult_125_B_not_8_port);
   mult_125_AN1_7_0 : inv port map( inb => input_sample_mem_7_port, outb => 
                           mult_125_B_not_7_port);
   mult_125_AN1_6_0 : inv port map( inb => input_sample_mem_6_port, outb => 
                           mult_125_B_not_6_port);
   mult_125_AN1_5_0 : inv port map( inb => input_sample_mem_5_port, outb => 
                           mult_125_B_not_5_port);
   mult_125_AN1_4_0 : inv port map( inb => input_sample_mem_4_port, outb => 
                           mult_125_B_not_4_port);
   mult_125_AN1_3_0 : inv port map( inb => input_sample_mem_3_port, outb => 
                           mult_125_B_not_3_port);
   mult_125_AN1_2_0 : inv port map( inb => input_sample_mem_2_port, outb => 
                           mult_125_B_not_2_port);
   mult_125_AN1_1_0 : inv port map( inb => input_sample_mem_1_port, outb => 
                           mult_125_B_not_1_port);
   mult_125_AN1_0_0 : inv port map( inb => input_sample_mem_0_port, outb => 
                           mult_125_B_not_0_port);
   mult_125_AN1_15_15 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_15_15_port);
   mult_125_AN3_15_14 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_14_port, outb => 
                           mult_125_ab_15_14_port);
   mult_125_AN3_15_13 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_13_port, outb => 
                           mult_125_ab_15_13_port);
   mult_125_AN3_15_12 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_12_port, outb => 
                           mult_125_ab_15_12_port);
   mult_125_AN3_15_11 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_11_port, outb => 
                           mult_125_ab_15_11_port);
   mult_125_AN3_15_10 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_10_port, outb => 
                           mult_125_ab_15_10_port);
   mult_125_AN3_15_9 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_9_port, outb => 
                           mult_125_ab_15_9_port);
   mult_125_AN3_15_8 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_8_port, outb => 
                           mult_125_ab_15_8_port);
   mult_125_AN3_15_7 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_7_port, outb => 
                           mult_125_ab_15_7_port);
   mult_125_AN3_15_6 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_6_port, outb => 
                           mult_125_ab_15_6_port);
   mult_125_AN3_15_5 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_5_port, outb => 
                           mult_125_ab_15_5_port);
   mult_125_AN3_15_4 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_4_port, outb => 
                           mult_125_ab_15_4_port);
   mult_125_AN3_15_3 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_3_port, outb => 
                           mult_125_ab_15_3_port);
   mult_125_AN3_15_2 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_2_port, outb => 
                           mult_125_ab_15_2_port);
   mult_125_AN3_15_1 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_1_port, outb => 
                           mult_125_ab_15_1_port);
   mult_125_AN3_15_0 : nor2 port map( a => mult_125_A_not_15_port, b => 
                           mult_125_B_notx_0_port, outb => 
                           mult_125_ab_15_0_port);
   mult_125_AN2_14_15 : nor2 port map( a => mult_125_A_notx_14_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_14_15_port);
   mult_125_AN1_14_14 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_14_14_port);
   mult_125_AN1_14_13 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_14_13_port);
   mult_125_AN1_14_12 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_14_12_port);
   mult_125_AN1_14_11 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_14_11_port);
   mult_125_AN1_14_10 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_14_10_port);
   mult_125_AN1_14_9 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_14_9_port
                           );
   mult_125_AN1_14_8 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_14_8_port
                           );
   mult_125_AN1_14_7 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_14_7_port
                           );
   mult_125_AN1_14_6 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_14_6_port
                           );
   mult_125_AN1_14_5 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_14_5_port
                           );
   mult_125_AN1_14_4 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_14_4_port
                           );
   mult_125_AN1_14_3 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_14_3_port
                           );
   mult_125_AN1_14_2 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_14_2_port
                           );
   mult_125_AN1_14_1 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_14_1_port
                           );
   mult_125_AN1_14_0_0 : nor2 port map( a => mult_125_A_not_14_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_14_0_port
                           );
   mult_125_AN2_13_15 : nor2 port map( a => mult_125_A_notx_13_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_13_15_port);
   mult_125_AN1_13_14 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_13_14_port);
   mult_125_AN1_13_13 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_13_13_port);
   mult_125_AN1_13_12 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_13_12_port);
   mult_125_AN1_13_11 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_13_11_port);
   mult_125_AN1_13_10 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_13_10_port);
   mult_125_AN1_13_9 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_13_9_port
                           );
   mult_125_AN1_13_8 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_13_8_port
                           );
   mult_125_AN1_13_7 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_13_7_port
                           );
   mult_125_AN1_13_6 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_13_6_port
                           );
   mult_125_AN1_13_5 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_13_5_port
                           );
   mult_125_AN1_13_4 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_13_4_port
                           );
   mult_125_AN1_13_3 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_13_3_port
                           );
   mult_125_AN1_13_2 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_13_2_port
                           );
   mult_125_AN1_13_1 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_13_1_port
                           );
   mult_125_AN1_13_0_0 : nor2 port map( a => mult_125_A_not_13_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_13_0_port
                           );
   mult_125_AN2_12_15 : nor2 port map( a => mult_125_A_notx_12_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_12_15_port);
   mult_125_AN1_12_14 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_12_14_port);
   mult_125_AN1_12_13 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_12_13_port);
   mult_125_AN1_12_12 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_12_12_port);
   mult_125_AN1_12_11 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_12_11_port);
   mult_125_AN1_12_10 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_12_10_port);
   mult_125_AN1_12_9 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_12_9_port
                           );
   mult_125_AN1_12_8 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_12_8_port
                           );
   mult_125_AN1_12_7 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_12_7_port
                           );
   mult_125_AN1_12_6 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_12_6_port
                           );
   mult_125_AN1_12_5 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_12_5_port
                           );
   mult_125_AN1_12_4 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_12_4_port
                           );
   mult_125_AN1_12_3 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_12_3_port
                           );
   mult_125_AN1_12_2 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_12_2_port
                           );
   mult_125_AN1_12_1 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_12_1_port
                           );
   mult_125_AN1_12_0_0 : nor2 port map( a => mult_125_A_not_12_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_12_0_port
                           );
   mult_125_AN2_11_15 : nor2 port map( a => mult_125_A_notx_11_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_11_15_port);
   mult_125_AN1_11_14 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_11_14_port);
   mult_125_AN1_11_13 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_11_13_port);
   mult_125_AN1_11_12 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_11_12_port);
   mult_125_AN1_11_11 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_11_11_port);
   mult_125_AN1_11_10 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_11_10_port);
   mult_125_AN1_11_9 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_11_9_port
                           );
   mult_125_AN1_11_8 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_11_8_port
                           );
   mult_125_AN1_11_7 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_11_7_port
                           );
   mult_125_AN1_11_6 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_11_6_port
                           );
   mult_125_AN1_11_5 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_11_5_port
                           );
   mult_125_AN1_11_4 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_11_4_port
                           );
   mult_125_AN1_11_3 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_11_3_port
                           );
   mult_125_AN1_11_2 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_11_2_port
                           );
   mult_125_AN1_11_1 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_11_1_port
                           );
   mult_125_AN1_11_0_0 : nor2 port map( a => mult_125_A_not_11_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_11_0_port
                           );
   mult_125_AN2_10_15 : nor2 port map( a => mult_125_A_notx_10_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_10_15_port);
   mult_125_AN1_10_14 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_10_14_port);
   mult_125_AN1_10_13 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_10_13_port);
   mult_125_AN1_10_12 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_10_12_port);
   mult_125_AN1_10_11 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_10_11_port);
   mult_125_AN1_10_10 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_10_10_port);
   mult_125_AN1_10_9 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_10_9_port
                           );
   mult_125_AN1_10_8 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_10_8_port
                           );
   mult_125_AN1_10_7 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_10_7_port
                           );
   mult_125_AN1_10_6 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_10_6_port
                           );
   mult_125_AN1_10_5 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_10_5_port
                           );
   mult_125_AN1_10_4 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_10_4_port
                           );
   mult_125_AN1_10_3 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_10_3_port
                           );
   mult_125_AN1_10_2 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_10_2_port
                           );
   mult_125_AN1_10_1 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_10_1_port
                           );
   mult_125_AN1_10_0_0 : nor2 port map( a => mult_125_A_not_10_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_10_0_port
                           );
   mult_125_AN2_9_15 : nor2 port map( a => mult_125_A_notx_9_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_9_15_port);
   mult_125_AN1_9_14 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_9_14_port);
   mult_125_AN1_9_13 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_9_13_port);
   mult_125_AN1_9_12 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_9_12_port);
   mult_125_AN1_9_11 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_9_11_port);
   mult_125_AN1_9_10 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_9_10_port);
   mult_125_AN1_9_9 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_9_9_port)
                           ;
   mult_125_AN1_9_8 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_9_8_port)
                           ;
   mult_125_AN1_9_7 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_9_7_port)
                           ;
   mult_125_AN1_9_6 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_9_6_port)
                           ;
   mult_125_AN1_9_5 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_9_5_port)
                           ;
   mult_125_AN1_9_4 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_9_4_port)
                           ;
   mult_125_AN1_9_3 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_9_3_port)
                           ;
   mult_125_AN1_9_2 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_9_2_port)
                           ;
   mult_125_AN1_9_1 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_9_1_port)
                           ;
   mult_125_AN1_9_0_0 : nor2 port map( a => mult_125_A_not_9_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_9_0_port)
                           ;
   mult_125_AN2_8_15 : nor2 port map( a => mult_125_A_notx_8_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_8_15_port);
   mult_125_AN1_8_14 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_8_14_port);
   mult_125_AN1_8_13 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_8_13_port);
   mult_125_AN1_8_12 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_8_12_port);
   mult_125_AN1_8_11 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_8_11_port);
   mult_125_AN1_8_10 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_8_10_port);
   mult_125_AN1_8_9 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_8_9_port)
                           ;
   mult_125_AN1_8_8 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_8_8_port)
                           ;
   mult_125_AN1_8_7 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_8_7_port)
                           ;
   mult_125_AN1_8_6 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_8_6_port)
                           ;
   mult_125_AN1_8_5 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_8_5_port)
                           ;
   mult_125_AN1_8_4 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_8_4_port)
                           ;
   mult_125_AN1_8_3 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_8_3_port)
                           ;
   mult_125_AN1_8_2 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_8_2_port)
                           ;
   mult_125_AN1_8_1 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_8_1_port)
                           ;
   mult_125_AN1_8_0_0 : nor2 port map( a => mult_125_A_not_8_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_8_0_port)
                           ;
   mult_125_AN2_7_15 : nor2 port map( a => mult_125_A_notx_7_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_7_15_port);
   mult_125_AN1_7_14 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_7_14_port);
   mult_125_AN1_7_13 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_7_13_port);
   mult_125_AN1_7_12 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_7_12_port);
   mult_125_AN1_7_11 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_7_11_port);
   mult_125_AN1_7_10 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_7_10_port);
   mult_125_AN1_7_9 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_7_9_port)
                           ;
   mult_125_AN1_7_8 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_7_8_port)
                           ;
   mult_125_AN1_7_7 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_7_7_port)
                           ;
   mult_125_AN1_7_6 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_7_6_port)
                           ;
   mult_125_AN1_7_5 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_7_5_port)
                           ;
   mult_125_AN1_7_4 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_7_4_port)
                           ;
   mult_125_AN1_7_3 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_7_3_port)
                           ;
   mult_125_AN1_7_2 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_7_2_port)
                           ;
   mult_125_AN1_7_1 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_7_1_port)
                           ;
   mult_125_AN1_7_0_0 : nor2 port map( a => mult_125_A_not_7_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_7_0_port)
                           ;
   mult_125_AN2_6_15 : nor2 port map( a => mult_125_A_notx_6_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_6_15_port);
   mult_125_AN1_6_14 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_6_14_port);
   mult_125_AN1_6_13 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_6_13_port);
   mult_125_AN1_6_12 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_6_12_port);
   mult_125_AN1_6_11 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_6_11_port);
   mult_125_AN1_6_10 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_6_10_port);
   mult_125_AN1_6_9 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_6_9_port)
                           ;
   mult_125_AN1_6_8 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_6_8_port)
                           ;
   mult_125_AN1_6_7 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_6_7_port)
                           ;
   mult_125_AN1_6_6 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_6_6_port)
                           ;
   mult_125_AN1_6_5 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_6_5_port)
                           ;
   mult_125_AN1_6_4 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_6_4_port)
                           ;
   mult_125_AN1_6_3 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_6_3_port)
                           ;
   mult_125_AN1_6_2 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_6_2_port)
                           ;
   mult_125_AN1_6_1 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_6_1_port)
                           ;
   mult_125_AN1_6_0_0 : nor2 port map( a => mult_125_A_not_6_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_6_0_port)
                           ;
   mult_125_AN2_5_15 : nor2 port map( a => mult_125_A_notx_5_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_5_15_port);
   mult_125_AN1_5_14 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_5_14_port);
   mult_125_AN1_5_13 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_5_13_port);
   mult_125_AN1_5_12 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_5_12_port);
   mult_125_AN1_5_11 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_5_11_port);
   mult_125_AN1_5_10 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_5_10_port);
   mult_125_AN1_5_9 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_5_9_port)
                           ;
   mult_125_AN1_5_8 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_5_8_port)
                           ;
   mult_125_AN1_5_7 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_5_7_port)
                           ;
   mult_125_AN1_5_6 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_5_6_port)
                           ;
   mult_125_AN1_5_5 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_5_5_port)
                           ;
   mult_125_AN1_5_4 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_5_4_port)
                           ;
   mult_125_AN1_5_3 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_5_3_port)
                           ;
   mult_125_AN1_5_2 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_5_2_port)
                           ;
   mult_125_AN1_5_1 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_5_1_port)
                           ;
   mult_125_AN1_5_0_0 : nor2 port map( a => mult_125_A_not_5_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_5_0_port)
                           ;
   mult_125_AN2_4_15 : nor2 port map( a => mult_125_A_notx_4_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_4_15_port);
   mult_125_AN1_4_14 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_4_14_port);
   mult_125_AN1_4_13 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_4_13_port);
   mult_125_AN1_4_12 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_4_12_port);
   mult_125_AN1_4_11 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_4_11_port);
   mult_125_AN1_4_10 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_4_10_port);
   mult_125_AN1_4_9 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_4_9_port)
                           ;
   mult_125_AN1_4_8 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_4_8_port)
                           ;
   mult_125_AN1_4_7 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_4_7_port)
                           ;
   mult_125_AN1_4_6 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_4_6_port)
                           ;
   mult_125_AN1_4_5 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_4_5_port)
                           ;
   mult_125_AN1_4_4 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_4_4_port)
                           ;
   mult_125_AN1_4_3 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_4_3_port)
                           ;
   mult_125_AN1_4_2 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_4_2_port)
                           ;
   mult_125_AN1_4_1 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_4_1_port)
                           ;
   mult_125_AN1_4_0_0 : nor2 port map( a => mult_125_A_not_4_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_4_0_port)
                           ;
   mult_125_AN2_3_15 : nor2 port map( a => mult_125_A_notx_3_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_3_15_port);
   mult_125_AN1_3_14 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_3_14_port);
   mult_125_AN1_3_13 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_3_13_port);
   mult_125_AN1_3_12 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_3_12_port);
   mult_125_AN1_3_11 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_3_11_port);
   mult_125_AN1_3_10 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_3_10_port);
   mult_125_AN1_3_9 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_3_9_port)
                           ;
   mult_125_AN1_3_8 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_3_8_port)
                           ;
   mult_125_AN1_3_7 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_3_7_port)
                           ;
   mult_125_AN1_3_6 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_3_6_port)
                           ;
   mult_125_AN1_3_5 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_3_5_port)
                           ;
   mult_125_AN1_3_4 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_3_4_port)
                           ;
   mult_125_AN1_3_3 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_3_3_port)
                           ;
   mult_125_AN1_3_2 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_3_2_port)
                           ;
   mult_125_AN1_3_1 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_3_1_port)
                           ;
   mult_125_AN1_3_0_0 : nor2 port map( a => mult_125_A_not_3_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_3_0_port)
                           ;
   mult_125_AN2_2_15 : nor2 port map( a => mult_125_A_notx_2_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_2_15_port);
   mult_125_AN1_2_14 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_2_14_port);
   mult_125_AN1_2_13 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_2_13_port);
   mult_125_AN1_2_12 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_2_12_port);
   mult_125_AN1_2_11 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_2_11_port);
   mult_125_AN1_2_10 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_2_10_port);
   mult_125_AN1_2_9 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_2_9_port)
                           ;
   mult_125_AN1_2_8 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_2_8_port)
                           ;
   mult_125_AN1_2_7 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_2_7_port)
                           ;
   mult_125_AN1_2_6 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_2_6_port)
                           ;
   mult_125_AN1_2_5 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_2_5_port)
                           ;
   mult_125_AN1_2_4 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_2_4_port)
                           ;
   mult_125_AN1_2_3 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_2_3_port)
                           ;
   mult_125_AN1_2_2 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_2_2_port)
                           ;
   mult_125_AN1_2_1 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_2_1_port)
                           ;
   mult_125_AN1_2_0_0 : nor2 port map( a => mult_125_A_not_2_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_2_0_port)
                           ;
   mult_125_AN2_1_15 : nor2 port map( a => mult_125_A_notx_1_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_1_15_port);
   mult_125_AN1_1_14 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_1_14_port);
   mult_125_AN1_1_13 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_1_13_port);
   mult_125_AN1_1_12 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_1_12_port);
   mult_125_AN1_1_11 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_1_11_port);
   mult_125_AN1_1_10 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_1_10_port);
   mult_125_AN1_1_9 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_1_9_port)
                           ;
   mult_125_AN1_1_8 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_1_8_port)
                           ;
   mult_125_AN1_1_7 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_1_7_port)
                           ;
   mult_125_AN1_1_6 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_1_6_port)
                           ;
   mult_125_AN1_1_5 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_1_5_port)
                           ;
   mult_125_AN1_1_4 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_1_4_port)
                           ;
   mult_125_AN1_1_3 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_1_3_port)
                           ;
   mult_125_AN1_1_2 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_1_2_port)
                           ;
   mult_125_AN1_1_1 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_1_1_port)
                           ;
   mult_125_AN1_1_0_0 : nor2 port map( a => mult_125_A_not_1_port, b => 
                           mult_125_B_not_0_port, outb => mult_125_ab_1_0_port)
                           ;
   mult_125_AN2_0_15 : nor2 port map( a => mult_125_A_notx_0_port, b => 
                           mult_125_B_not_15_port, outb => 
                           mult_125_ab_0_15_port);
   mult_125_AN1_0_14 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_14_port, outb => 
                           mult_125_ab_0_14_port);
   mult_125_AN1_0_13 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_13_port, outb => 
                           mult_125_ab_0_13_port);
   mult_125_AN1_0_12 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_12_port, outb => 
                           mult_125_ab_0_12_port);
   mult_125_AN1_0_11 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_11_port, outb => 
                           mult_125_ab_0_11_port);
   mult_125_AN1_0_10 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_10_port, outb => 
                           mult_125_ab_0_10_port);
   mult_125_AN1_0_9 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_9_port, outb => mult_125_ab_0_9_port)
                           ;
   mult_125_AN1_0_8 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_8_port, outb => mult_125_ab_0_8_port)
                           ;
   mult_125_AN1_0_7 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_7_port, outb => mult_125_ab_0_7_port)
                           ;
   mult_125_AN1_0_6 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_6_port, outb => mult_125_ab_0_6_port)
                           ;
   mult_125_AN1_0_5 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_5_port, outb => mult_125_ab_0_5_port)
                           ;
   mult_125_AN1_0_4 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_4_port, outb => mult_125_ab_0_4_port)
                           ;
   mult_125_AN1_0_3 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_3_port, outb => mult_125_ab_0_3_port)
                           ;
   mult_125_AN1_0_2 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_2_port, outb => mult_125_ab_0_2_port)
                           ;
   mult_125_AN1_0_1 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_1_port, outb => mult_125_ab_0_1_port)
                           ;
   mult_125_AN1_0_0_0 : nor2 port map( a => mult_125_A_not_0_port, b => 
                           mult_125_B_not_0_port, outb => 
                           multiplier_sigs_0_0_port);
   mult_125_G4_FS_1_U6_1_1_3 : oai12 port map( b => n5657, c => n5658, a => 
                           n5659, outb => mult_125_G4_FS_1_C_1_7_0_port);
   mult_125_G4_FS_1_U6_1_1_2 : oai12 port map( b => n5654, c => n5655, a => 
                           n5656, outb => mult_125_G4_FS_1_C_1_6_0_port);
   mult_125_G4_FS_1_U6_1_1_1 : oai12 port map( b => n5651, c => n5652, a => 
                           n5653, outb => mult_125_G4_FS_1_C_1_5_0_port);
   mult_125_G4_FS_1_U6_0_7_1 : oai12 port map( b => n5648, c => n5649, a => 
                           mult_125_G4_FS_1_G_n_int_0_7_0_port, outb => 
                           mult_125_G4_FS_1_C_1_7_1_port);
   mult_125_G4_FS_1_U3_C_0_7_1 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_7_1_port, b => 
                           mult_125_G4_FS_1_C_1_7_1_port, outb => 
                           multiplier_sigs_3_31_port);
   mult_125_G4_FS_1_U3_B_0_7_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_7_1_port, b => 
                           mult_125_G4_FS_1_P_0_7_1_port, outb => n5647);
   mult_125_G4_FS_1_U2_0_7_1 : nand2 port map( a => mult_125_G4_A1_29_port, b 
                           => mult_125_G4_A2_29_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_7_1_port);
   mult_125_G4_FS_1_U1_0_7_1 : nand2 port map( a => n5645, b => n5646, outb => 
                           mult_125_G4_FS_1_P_0_7_1_port);
   mult_125_G4_FS_1_U3_C_0_7_0 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_7_0_port, b => 
                           mult_125_G4_FS_1_C_1_7_0_port, outb => 
                           multiplier_sigs_3_30_port);
   mult_125_G4_FS_1_U3_B_0_7_0 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_7_0_port, b => 
                           mult_125_G4_FS_1_TEMP_P_0_7_0_port, outb => n5644);
   mult_125_G4_FS_1_U2_0_7_0 : nand2 port map( a => mult_125_G4_A1_28_port, b 
                           => mult_125_G4_A2_28_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_7_0_port);
   mult_125_G4_FS_1_U1_0_7_0 : nand2 port map( a => n5642, b => n5643, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_7_0_port);
   mult_125_G4_FS_1_U6_0_6_3 : oai12 port map( b => n5640, c => n5641, a => 
                           mult_125_G4_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G4_FS_1_C_1_6_3_port);
   mult_125_G4_FS_1_U5_0_6_3 : oai12 port map( b => n5638, c => n5639, a => 
                           mult_125_G4_FS_1_G_n_int_0_6_3_port, outb => 
                           mult_125_G4_FS_1_G_1_1_2_port);
   mult_125_G4_FS_1_U4_0_6_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_6_2_port, b => 
                           mult_125_G4_FS_1_P_0_6_3_port, outb => n5658);
   mult_125_G4_FS_1_U3_C_0_6_3 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_6_3_port, b => 
                           mult_125_G4_FS_1_C_1_6_3_port, outb => 
                           multiplier_sigs_3_29_port);
   mult_125_G4_FS_1_U3_B_0_6_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_6_3_port, b => 
                           mult_125_G4_FS_1_P_0_6_3_port, outb => n5637);
   mult_125_G4_FS_1_U2_0_6_3 : nand2 port map( a => mult_125_G4_A1_27_port, b 
                           => mult_125_G4_A2_27_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_6_3_port);
   mult_125_G4_FS_1_U1_0_6_3 : nand2 port map( a => n5635, b => n5636, outb => 
                           mult_125_G4_FS_1_P_0_6_3_port);
   mult_125_G4_FS_1_U6_0_6_2 : oai12 port map( b => n5633, c => n5634, a => 
                           mult_125_G4_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G4_FS_1_C_1_6_2_port);
   mult_125_G4_FS_1_U5_0_6_2 : oai12 port map( b => n5632, c => n5641, a => 
                           mult_125_G4_FS_1_G_n_int_0_6_2_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_6_2_port);
   mult_125_G4_FS_1_U4_0_6_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_6_1_port, b => 
                           mult_125_G4_FS_1_P_0_6_2_port, outb => n5631);
   mult_125_G4_FS_1_U3_C_0_6_2 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_6_2_port, b => 
                           mult_125_G4_FS_1_C_1_6_2_port, outb => 
                           multiplier_sigs_3_28_port);
   mult_125_G4_FS_1_U3_B_0_6_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_6_2_port, b => 
                           mult_125_G4_FS_1_P_0_6_2_port, outb => n5630);
   mult_125_G4_FS_1_U2_0_6_2 : nand2 port map( a => mult_125_G4_A1_26_port, b 
                           => mult_125_G4_A2_26_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_6_2_port);
   mult_125_G4_FS_1_U1_0_6_2 : nand2 port map( a => n5628, b => n5629, outb => 
                           mult_125_G4_FS_1_P_0_6_2_port);
   mult_125_G4_FS_1_U6_0_6_1 : oai12 port map( b => n5657, c => n5627, a => 
                           mult_125_G4_FS_1_G_n_int_0_6_0_port, outb => 
                           mult_125_G4_FS_1_C_1_6_1_port);
   mult_125_G4_FS_1_U5_0_6_1 : oai12 port map( b => 
                           mult_125_G4_FS_1_G_n_int_0_6_0_port, c => n5634, a 
                           => mult_125_G4_FS_1_G_n_int_0_6_1_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_6_1_port);
   mult_125_G4_FS_1_U4_0_6_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_6_0_port, b => 
                           mult_125_G4_FS_1_P_0_6_1_port, outb => n5626);
   mult_125_G4_FS_1_U3_C_0_6_1 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_6_1_port, b => 
                           mult_125_G4_FS_1_C_1_6_1_port, outb => 
                           multiplier_sigs_3_27_port);
   mult_125_G4_FS_1_U3_B_0_6_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_6_1_port, b => 
                           mult_125_G4_FS_1_P_0_6_1_port, outb => n5625);
   mult_125_G4_FS_1_U2_0_6_1 : nand2 port map( a => mult_125_G4_A1_25_port, b 
                           => mult_125_G4_A2_25_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_6_1_port);
   mult_125_G4_FS_1_U1_0_6_1 : nand2 port map( a => n5623, b => n5624, outb => 
                           mult_125_G4_FS_1_P_0_6_1_port);
   mult_125_G4_FS_1_U3_C_0_6_0 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_6_0_port, b => 
                           mult_125_G4_FS_1_C_1_6_0_port, outb => 
                           multiplier_sigs_3_26_port);
   mult_125_G4_FS_1_U3_B_0_6_0 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_6_0_port, b => 
                           mult_125_G4_FS_1_TEMP_P_0_6_0_port, outb => n5622);
   mult_125_G4_FS_1_U2_0_6_0 : nand2 port map( a => mult_125_G4_A1_24_port, b 
                           => mult_125_G4_A2_24_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_6_0_port);
   mult_125_G4_FS_1_U1_0_6_0 : nand2 port map( a => n5620, b => n5621, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_6_0_port);
   mult_125_G4_FS_1_U6_0_5_3 : oai12 port map( b => n5618, c => n5619, a => 
                           mult_125_G4_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G4_FS_1_C_1_5_3_port);
   mult_125_G4_FS_1_U5_0_5_3 : oai12 port map( b => n5616, c => n5617, a => 
                           mult_125_G4_FS_1_G_n_int_0_5_3_port, outb => 
                           mult_125_G4_FS_1_G_1_1_1_port);
   mult_125_G4_FS_1_U4_0_5_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_5_2_port, b => 
                           mult_125_G4_FS_1_P_0_5_3_port, outb => n5655);
   mult_125_G4_FS_1_U3_C_0_5_3 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_5_3_port, b => 
                           mult_125_G4_FS_1_C_1_5_3_port, outb => 
                           multiplier_sigs_3_25_port);
   mult_125_G4_FS_1_U3_B_0_5_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_5_3_port, b => 
                           mult_125_G4_FS_1_P_0_5_3_port, outb => n5615);
   mult_125_G4_FS_1_U2_0_5_3 : nand2 port map( a => mult_125_G4_A1_23_port, b 
                           => mult_125_G4_A2_23_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_5_3_port);
   mult_125_G4_FS_1_U1_0_5_3 : nand2 port map( a => n5613, b => n5614, outb => 
                           mult_125_G4_FS_1_P_0_5_3_port);
   mult_125_G4_FS_1_U6_0_5_2 : oai12 port map( b => n5611, c => n5612, a => 
                           mult_125_G4_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G4_FS_1_C_1_5_2_port);
   mult_125_G4_FS_1_U5_0_5_2 : oai12 port map( b => n5610, c => n5619, a => 
                           mult_125_G4_FS_1_G_n_int_0_5_2_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_5_2_port);
   mult_125_G4_FS_1_U4_0_5_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_5_1_port, b => 
                           mult_125_G4_FS_1_P_0_5_2_port, outb => n5609);
   mult_125_G4_FS_1_U3_C_0_5_2 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_5_2_port, b => 
                           mult_125_G4_FS_1_C_1_5_2_port, outb => 
                           multiplier_sigs_3_24_port);
   mult_125_G4_FS_1_U3_B_0_5_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_5_2_port, b => 
                           mult_125_G4_FS_1_P_0_5_2_port, outb => n5608);
   mult_125_G4_FS_1_U2_0_5_2 : nand2 port map( a => mult_125_G4_A1_22_port, b 
                           => mult_125_G4_A2_22_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_5_2_port);
   mult_125_G4_FS_1_U1_0_5_2 : nand2 port map( a => n5606, b => n5607, outb => 
                           mult_125_G4_FS_1_P_0_5_2_port);
   mult_125_G4_FS_1_U6_0_5_1 : oai12 port map( b => n5654, c => n5605, a => 
                           mult_125_G4_FS_1_G_n_int_0_5_0_port, outb => 
                           mult_125_G4_FS_1_C_1_5_1_port);
   mult_125_G4_FS_1_U5_0_5_1 : oai12 port map( b => 
                           mult_125_G4_FS_1_G_n_int_0_5_0_port, c => n5612, a 
                           => mult_125_G4_FS_1_G_n_int_0_5_1_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_5_1_port);
   mult_125_G4_FS_1_U4_0_5_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_5_0_port, b => 
                           mult_125_G4_FS_1_P_0_5_1_port, outb => n5604);
   mult_125_G4_FS_1_U3_C_0_5_1 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_5_1_port, b => 
                           mult_125_G4_FS_1_C_1_5_1_port, outb => 
                           multiplier_sigs_3_23_port);
   mult_125_G4_FS_1_U3_B_0_5_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_5_1_port, b => 
                           mult_125_G4_FS_1_P_0_5_1_port, outb => n5603);
   mult_125_G4_FS_1_U2_0_5_1 : nand2 port map( a => mult_125_G4_A1_21_port, b 
                           => mult_125_G4_A2_21_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_5_1_port);
   mult_125_G4_FS_1_U1_0_5_1 : nand2 port map( a => n5601, b => n5602, outb => 
                           mult_125_G4_FS_1_P_0_5_1_port);
   mult_125_G4_FS_1_U3_C_0_5_0 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_5_0_port, b => 
                           mult_125_G4_FS_1_C_1_5_0_port, outb => 
                           multiplier_sigs_3_22_port);
   mult_125_G4_FS_1_U3_B_0_5_0 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_5_0_port, b => 
                           mult_125_G4_FS_1_TEMP_P_0_5_0_port, outb => n5600);
   mult_125_G4_FS_1_U2_0_5_0 : nand2 port map( a => mult_125_G4_A1_20_port, b 
                           => mult_125_G4_A2_20_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_5_0_port);
   mult_125_G4_FS_1_U1_0_5_0 : nand2 port map( a => n5598, b => n5599, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_5_0_port);
   mult_125_G4_FS_1_U6_0_4_3 : oai12 port map( b => n5596, c => n5597, a => 
                           mult_125_G4_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G4_FS_1_C_1_4_3_port);
   mult_125_G4_FS_1_U5_0_4_3 : oai12 port map( b => n5594, c => n5595, a => 
                           mult_125_G4_FS_1_G_n_int_0_4_3_port, outb => 
                           mult_125_G4_FS_1_G_1_1_0_port);
   mult_125_G4_FS_1_U4_0_4_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_4_2_port, b => 
                           mult_125_G4_FS_1_P_0_4_3_port, outb => n5652);
   mult_125_G4_FS_1_U3_C_0_4_3 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_4_3_port, b => 
                           mult_125_G4_FS_1_C_1_4_3_port, outb => 
                           multiplier_sigs_3_21_port);
   mult_125_G4_FS_1_U3_B_0_4_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_4_3_port, b => 
                           mult_125_G4_FS_1_P_0_4_3_port, outb => n5593);
   mult_125_G4_FS_1_U2_0_4_3 : nand2 port map( a => mult_125_G4_A1_19_port, b 
                           => mult_125_G4_A2_19_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_4_3_port);
   mult_125_G4_FS_1_U1_0_4_3 : nand2 port map( a => n5591, b => n5592, outb => 
                           mult_125_G4_FS_1_P_0_4_3_port);
   mult_125_G4_FS_1_U6_0_4_2 : oai12 port map( b => n5589, c => n5590, a => 
                           mult_125_G4_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G4_FS_1_C_1_4_2_port);
   mult_125_G4_FS_1_U5_0_4_2 : oai12 port map( b => n5588, c => n5597, a => 
                           mult_125_G4_FS_1_G_n_int_0_4_2_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_4_2_port);
   mult_125_G4_FS_1_U4_0_4_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_4_1_port, b => 
                           mult_125_G4_FS_1_P_0_4_2_port, outb => n5587);
   mult_125_G4_FS_1_U3_C_0_4_2 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_4_2_port, b => 
                           mult_125_G4_FS_1_C_1_4_2_port, outb => 
                           multiplier_sigs_3_20_port);
   mult_125_G4_FS_1_U3_B_0_4_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_4_2_port, b => 
                           mult_125_G4_FS_1_P_0_4_2_port, outb => n5586);
   mult_125_G4_FS_1_U2_0_4_2 : nand2 port map( a => mult_125_G4_A1_18_port, b 
                           => mult_125_G4_A2_18_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_4_2_port);
   mult_125_G4_FS_1_U1_0_4_2 : nand2 port map( a => n5584, b => n5585, outb => 
                           mult_125_G4_FS_1_P_0_4_2_port);
   mult_125_G4_FS_1_U6_0_4_1 : oai12 port map( b => n5651, c => n5583, a => 
                           mult_125_G4_FS_1_G_n_int_0_4_0_port, outb => 
                           mult_125_G4_FS_1_C_1_4_1_port);
   mult_125_G4_FS_1_U5_0_4_1 : oai12 port map( b => 
                           mult_125_G4_FS_1_G_n_int_0_4_0_port, c => n5590, a 
                           => mult_125_G4_FS_1_G_n_int_0_4_1_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_4_1_port);
   mult_125_G4_FS_1_U4_0_4_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_TEMP_P_0_4_0_port, b => 
                           mult_125_G4_FS_1_P_0_4_1_port, outb => n5582);
   mult_125_G4_FS_1_U3_C_0_4_1 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_4_1_port, b => 
                           mult_125_G4_FS_1_C_1_4_1_port, outb => 
                           multiplier_sigs_3_19_port);
   mult_125_G4_FS_1_U3_B_0_4_1 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_4_1_port, b => 
                           mult_125_G4_FS_1_P_0_4_1_port, outb => n5581);
   mult_125_G4_FS_1_U2_0_4_1 : nand2 port map( a => mult_125_G4_A1_17_port, b 
                           => mult_125_G4_A2_17_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_4_1_port);
   mult_125_G4_FS_1_U1_0_4_1 : nand2 port map( a => n5579, b => n5580, outb => 
                           mult_125_G4_FS_1_P_0_4_1_port);
   mult_125_G4_FS_1_U3_C_0_4_0 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_4_0_port, b => 
                           mult_125_G4_FS_1_C_1_4_0_port, outb => 
                           multiplier_sigs_3_18_port);
   mult_125_G4_FS_1_U3_B_0_4_0 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_4_0_port, b => 
                           mult_125_G4_FS_1_TEMP_P_0_4_0_port, outb => n5578);
   mult_125_G4_FS_1_U2_0_4_0 : nand2 port map( a => mult_125_G4_A1_16_port, b 
                           => mult_125_G4_A2_16_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_4_0_port);
   mult_125_G4_FS_1_U1_0_4_0 : nand2 port map( a => n5576, b => n5577, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_4_0_port);
   mult_125_G4_FS_1_U5_0_3_3 : oai12 port map( b => n5574, c => n5575, a => 
                           mult_125_G4_FS_1_G_n_int_0_3_3_port, outb => 
                           mult_125_G4_FS_1_G_1_0_3_port);
   mult_125_G4_FS_1_U3_C_0_3_3 : xor2 port map( a => 
                           mult_125_G4_FS_1_PG_int_0_3_3_port, b => 
                           mult_125_G4_FS_1_C_1_3_3_port, outb => 
                           multiplier_sigs_3_17_port);
   mult_125_G4_FS_1_U3_B_0_3_3 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_3_3_port, b => 
                           mult_125_G4_FS_1_P_0_3_3_port, outb => n5573);
   mult_125_G4_FS_1_U2_0_3_3 : nand2 port map( a => mult_125_G4_A1_15_port, b 
                           => mult_125_G4_A2_15_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_3_3_port);
   mult_125_G4_FS_1_U1_0_3_3 : nand2 port map( a => n5571, b => n5572, outb => 
                           mult_125_G4_FS_1_P_0_3_3_port);
   mult_125_G4_FS_1_U3_B_0_3_2 : nand2 port map( a => 
                           mult_125_G4_FS_1_G_n_int_0_3_2_port, b => 
                           mult_125_G4_FS_1_P_0_3_2_port, outb => n5570);
   mult_125_G4_FS_1_U2_0_3_2 : nand2 port map( a => mult_125_G4_A1_14_port, b 
                           => mult_125_G4_A2_14_port, outb => 
                           mult_125_G4_FS_1_G_n_int_0_3_2_port);
   mult_125_G4_FS_1_U1_0_3_2 : nand2 port map( a => n5568, b => n5569, outb => 
                           mult_125_G4_FS_1_P_0_3_2_port);
   mult_125_G4_AN1_15 : inv port map( inb => coefficient_mem_array_3_15_port, 
                           outb => mult_125_G4_A_not_15_port);
   mult_125_G4_AN1_14 : inv port map( inb => coefficient_mem_array_3_14_port, 
                           outb => mult_125_G4_A_not_14_port);
   mult_125_G4_AN1_13 : inv port map( inb => coefficient_mem_array_3_13_port, 
                           outb => mult_125_G4_A_not_13_port);
   mult_125_G4_AN1_12 : inv port map( inb => coefficient_mem_array_3_12_port, 
                           outb => mult_125_G4_A_not_12_port);
   mult_125_G4_AN1_11 : inv port map( inb => coefficient_mem_array_3_11_port, 
                           outb => mult_125_G4_A_not_11_port);
   mult_125_G4_AN1_10 : inv port map( inb => coefficient_mem_array_3_10_port, 
                           outb => mult_125_G4_A_not_10_port);
   mult_125_G4_AN1_9 : inv port map( inb => coefficient_mem_array_3_9_port, 
                           outb => mult_125_G4_A_not_9_port);
   mult_125_G4_AN1_8 : inv port map( inb => coefficient_mem_array_3_8_port, 
                           outb => mult_125_G4_A_not_8_port);
   mult_125_G4_AN1_7 : inv port map( inb => coefficient_mem_array_3_7_port, 
                           outb => mult_125_G4_A_not_7_port);
   mult_125_G4_AN1_6 : inv port map( inb => coefficient_mem_array_3_6_port, 
                           outb => mult_125_G4_A_not_6_port);
   mult_125_G4_AN1_5 : inv port map( inb => coefficient_mem_array_3_5_port, 
                           outb => mult_125_G4_A_not_5_port);
   mult_125_G4_AN1_4 : inv port map( inb => coefficient_mem_array_3_4_port, 
                           outb => mult_125_G4_A_not_4_port);
   mult_125_G4_AN1_3 : inv port map( inb => coefficient_mem_array_3_3_port, 
                           outb => mult_125_G4_A_not_3_port);
   mult_125_G4_AN1_2 : inv port map( inb => coefficient_mem_array_3_2_port, 
                           outb => mult_125_G4_A_not_2_port);
   mult_125_G4_AN1_1 : inv port map( inb => coefficient_mem_array_3_1_port, 
                           outb => mult_125_G4_A_not_1_port);
   mult_125_G4_AN1_0 : inv port map( inb => coefficient_mem_array_3_0_port, 
                           outb => mult_125_G4_A_not_0_port);
   mult_125_G4_AN1_15_0 : inv port map( inb => input_sample_mem_15_port, outb 
                           => mult_125_G4_B_not_15_port);
   mult_125_G4_AN1_14_0 : inv port map( inb => input_sample_mem_14_port, outb 
                           => mult_125_G4_B_not_14_port);
   mult_125_G4_AN1_13_0 : inv port map( inb => input_sample_mem_13_port, outb 
                           => mult_125_G4_B_not_13_port);
   mult_125_G4_AN1_12_0 : inv port map( inb => input_sample_mem_12_port, outb 
                           => mult_125_G4_B_not_12_port);
   mult_125_G4_AN1_11_0 : inv port map( inb => input_sample_mem_11_port, outb 
                           => mult_125_G4_B_not_11_port);
   mult_125_G4_AN1_10_0 : inv port map( inb => input_sample_mem_10_port, outb 
                           => mult_125_G4_B_not_10_port);
   mult_125_G4_AN1_9_0 : inv port map( inb => input_sample_mem_9_port, outb => 
                           mult_125_G4_B_not_9_port);
   mult_125_G4_AN1_8_0 : inv port map( inb => input_sample_mem_8_port, outb => 
                           mult_125_G4_B_not_8_port);
   mult_125_G4_AN1_7_0 : inv port map( inb => input_sample_mem_7_port, outb => 
                           mult_125_G4_B_not_7_port);
   mult_125_G4_AN1_6_0 : inv port map( inb => input_sample_mem_6_port, outb => 
                           mult_125_G4_B_not_6_port);
   mult_125_G4_AN1_5_0 : inv port map( inb => input_sample_mem_5_port, outb => 
                           mult_125_G4_B_not_5_port);
   mult_125_G4_AN1_4_0 : inv port map( inb => input_sample_mem_4_port, outb => 
                           mult_125_G4_B_not_4_port);
   mult_125_G4_AN1_3_0 : inv port map( inb => input_sample_mem_3_port, outb => 
                           mult_125_G4_B_not_3_port);
   mult_125_G4_AN1_2_0 : inv port map( inb => input_sample_mem_2_port, outb => 
                           mult_125_G4_B_not_2_port);
   mult_125_G4_AN1_1_0 : inv port map( inb => input_sample_mem_1_port, outb => 
                           mult_125_G4_B_not_1_port);
   mult_125_G4_AN1_0_0 : inv port map( inb => input_sample_mem_0_port, outb => 
                           mult_125_G4_B_not_0_port);
   mult_125_G4_AN1_15_15 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_15_15_port);
   mult_125_G4_AN3_15_14 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_14_port, outb => 
                           mult_125_G4_ab_15_14_port);
   mult_125_G4_AN3_15_13 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_13_port, outb => 
                           mult_125_G4_ab_15_13_port);
   mult_125_G4_AN3_15_12 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_12_port, outb => 
                           mult_125_G4_ab_15_12_port);
   mult_125_G4_AN3_15_11 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_11_port, outb => 
                           mult_125_G4_ab_15_11_port);
   mult_125_G4_AN3_15_10 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_10_port, outb => 
                           mult_125_G4_ab_15_10_port);
   mult_125_G4_AN3_15_9 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_9_port, outb => 
                           mult_125_G4_ab_15_9_port);
   mult_125_G4_AN3_15_8 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_8_port, outb => 
                           mult_125_G4_ab_15_8_port);
   mult_125_G4_AN3_15_7 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_7_port, outb => 
                           mult_125_G4_ab_15_7_port);
   mult_125_G4_AN3_15_6 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_6_port, outb => 
                           mult_125_G4_ab_15_6_port);
   mult_125_G4_AN3_15_5 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_5_port, outb => 
                           mult_125_G4_ab_15_5_port);
   mult_125_G4_AN3_15_4 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_4_port, outb => 
                           mult_125_G4_ab_15_4_port);
   mult_125_G4_AN3_15_3 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_3_port, outb => 
                           mult_125_G4_ab_15_3_port);
   mult_125_G4_AN3_15_2 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_2_port, outb => 
                           mult_125_G4_ab_15_2_port);
   mult_125_G4_AN3_15_1 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_1_port, outb => 
                           mult_125_G4_ab_15_1_port);
   mult_125_G4_AN3_15_0 : nor2 port map( a => mult_125_G4_A_not_15_port, b => 
                           mult_125_G4_B_notx_0_port, outb => 
                           mult_125_G4_ab_15_0_port);
   mult_125_G4_AN2_14_15 : nor2 port map( a => mult_125_G4_A_notx_14_port, b =>
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_14_15_port);
   mult_125_G4_AN1_14_14 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_14_14_port);
   mult_125_G4_AN1_14_13 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_14_13_port);
   mult_125_G4_AN1_14_12 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_14_12_port);
   mult_125_G4_AN1_14_11 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_14_11_port);
   mult_125_G4_AN1_14_10 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_14_10_port);
   mult_125_G4_AN1_14_9 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_14_9_port);
   mult_125_G4_AN1_14_8 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_14_8_port);
   mult_125_G4_AN1_14_7 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_14_7_port);
   mult_125_G4_AN1_14_6 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_14_6_port);
   mult_125_G4_AN1_14_5 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_14_5_port);
   mult_125_G4_AN1_14_4 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_14_4_port);
   mult_125_G4_AN1_14_3 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_14_3_port);
   mult_125_G4_AN1_14_2 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_14_2_port);
   mult_125_G4_AN1_14_1 : nor2 port map( a => mult_125_G4_A_not_14_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_14_1_port);
   mult_125_G4_AN1_14_0_0 : nor2 port map( a => mult_125_G4_A_not_14_port, b =>
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_14_0_port);
   mult_125_G4_AN2_13_15 : nor2 port map( a => mult_125_G4_A_notx_13_port, b =>
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_13_15_port);
   mult_125_G4_AN1_13_14 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_13_14_port);
   mult_125_G4_AN1_13_13 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_13_13_port);
   mult_125_G4_AN1_13_12 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_13_12_port);
   mult_125_G4_AN1_13_11 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_13_11_port);
   mult_125_G4_AN1_13_10 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_13_10_port);
   mult_125_G4_AN1_13_9 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_13_9_port);
   mult_125_G4_AN1_13_8 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_13_8_port);
   mult_125_G4_AN1_13_7 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_13_7_port);
   mult_125_G4_AN1_13_6 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_13_6_port);
   mult_125_G4_AN1_13_5 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_13_5_port);
   mult_125_G4_AN1_13_4 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_13_4_port);
   mult_125_G4_AN1_13_3 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_13_3_port);
   mult_125_G4_AN1_13_2 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_13_2_port);
   mult_125_G4_AN1_13_1 : nor2 port map( a => mult_125_G4_A_not_13_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_13_1_port);
   mult_125_G4_AN1_13_0_0 : nor2 port map( a => mult_125_G4_A_not_13_port, b =>
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_13_0_port);
   mult_125_G4_AN2_12_15 : nor2 port map( a => mult_125_G4_A_notx_12_port, b =>
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_12_15_port);
   mult_125_G4_AN1_12_14 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_12_14_port);
   mult_125_G4_AN1_12_13 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_12_13_port);
   mult_125_G4_AN1_12_12 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_12_12_port);
   mult_125_G4_AN1_12_11 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_12_11_port);
   mult_125_G4_AN1_12_10 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_12_10_port);
   mult_125_G4_AN1_12_9 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_12_9_port);
   mult_125_G4_AN1_12_8 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_12_8_port);
   mult_125_G4_AN1_12_7 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_12_7_port);
   mult_125_G4_AN1_12_6 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_12_6_port);
   mult_125_G4_AN1_12_5 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_12_5_port);
   mult_125_G4_AN1_12_4 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_12_4_port);
   mult_125_G4_AN1_12_3 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_12_3_port);
   mult_125_G4_AN1_12_2 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_12_2_port);
   mult_125_G4_AN1_12_1 : nor2 port map( a => mult_125_G4_A_not_12_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_12_1_port);
   mult_125_G4_AN1_12_0_0 : nor2 port map( a => mult_125_G4_A_not_12_port, b =>
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_12_0_port);
   mult_125_G4_AN2_11_15 : nor2 port map( a => mult_125_G4_A_notx_11_port, b =>
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_11_15_port);
   mult_125_G4_AN1_11_14 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_11_14_port);
   mult_125_G4_AN1_11_13 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_11_13_port);
   mult_125_G4_AN1_11_12 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_11_12_port);
   mult_125_G4_AN1_11_11 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_11_11_port);
   mult_125_G4_AN1_11_10 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_11_10_port);
   mult_125_G4_AN1_11_9 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_11_9_port);
   mult_125_G4_AN1_11_8 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_11_8_port);
   mult_125_G4_AN1_11_7 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_11_7_port);
   mult_125_G4_AN1_11_6 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_11_6_port);
   mult_125_G4_AN1_11_5 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_11_5_port);
   mult_125_G4_AN1_11_4 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_11_4_port);
   mult_125_G4_AN1_11_3 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_11_3_port);
   mult_125_G4_AN1_11_2 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_11_2_port);
   mult_125_G4_AN1_11_1 : nor2 port map( a => mult_125_G4_A_not_11_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_11_1_port);
   mult_125_G4_AN1_11_0_0 : nor2 port map( a => mult_125_G4_A_not_11_port, b =>
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_11_0_port);
   mult_125_G4_AN2_10_15 : nor2 port map( a => mult_125_G4_A_notx_10_port, b =>
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_10_15_port);
   mult_125_G4_AN1_10_14 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_10_14_port);
   mult_125_G4_AN1_10_13 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_10_13_port);
   mult_125_G4_AN1_10_12 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_10_12_port);
   mult_125_G4_AN1_10_11 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_10_11_port);
   mult_125_G4_AN1_10_10 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_10_10_port);
   mult_125_G4_AN1_10_9 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_10_9_port);
   mult_125_G4_AN1_10_8 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_10_8_port);
   mult_125_G4_AN1_10_7 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_10_7_port);
   mult_125_G4_AN1_10_6 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_10_6_port);
   mult_125_G4_AN1_10_5 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_10_5_port);
   mult_125_G4_AN1_10_4 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_10_4_port);
   mult_125_G4_AN1_10_3 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_10_3_port);
   mult_125_G4_AN1_10_2 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_10_2_port);
   mult_125_G4_AN1_10_1 : nor2 port map( a => mult_125_G4_A_not_10_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_10_1_port);
   mult_125_G4_AN1_10_0_0 : nor2 port map( a => mult_125_G4_A_not_10_port, b =>
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_10_0_port);
   mult_125_G4_AN2_9_15 : nor2 port map( a => mult_125_G4_A_notx_9_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_9_15_port);
   mult_125_G4_AN1_9_14 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_9_14_port);
   mult_125_G4_AN1_9_13 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_9_13_port);
   mult_125_G4_AN1_9_12 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_9_12_port);
   mult_125_G4_AN1_9_11 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_9_11_port);
   mult_125_G4_AN1_9_10 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_9_10_port);
   mult_125_G4_AN1_9_9 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_9_9_port);
   mult_125_G4_AN1_9_8 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_9_8_port);
   mult_125_G4_AN1_9_7 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_9_7_port);
   mult_125_G4_AN1_9_6 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_9_6_port);
   mult_125_G4_AN1_9_5 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_9_5_port);
   mult_125_G4_AN1_9_4 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_9_4_port);
   mult_125_G4_AN1_9_3 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_9_3_port);
   mult_125_G4_AN1_9_2 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_9_2_port);
   mult_125_G4_AN1_9_1 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_9_1_port);
   mult_125_G4_AN1_9_0_0 : nor2 port map( a => mult_125_G4_A_not_9_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_9_0_port);
   mult_125_G4_AN2_8_15 : nor2 port map( a => mult_125_G4_A_notx_8_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_8_15_port);
   mult_125_G4_AN1_8_14 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_8_14_port);
   mult_125_G4_AN1_8_13 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_8_13_port);
   mult_125_G4_AN1_8_12 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_8_12_port);
   mult_125_G4_AN1_8_11 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_8_11_port);
   mult_125_G4_AN1_8_10 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_8_10_port);
   mult_125_G4_AN1_8_9 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_8_9_port);
   mult_125_G4_AN1_8_8 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_8_8_port);
   mult_125_G4_AN1_8_7 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_8_7_port);
   mult_125_G4_AN1_8_6 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_8_6_port);
   mult_125_G4_AN1_8_5 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_8_5_port);
   mult_125_G4_AN1_8_4 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_8_4_port);
   mult_125_G4_AN1_8_3 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_8_3_port);
   mult_125_G4_AN1_8_2 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_8_2_port);
   mult_125_G4_AN1_8_1 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_8_1_port);
   mult_125_G4_AN1_8_0_0 : nor2 port map( a => mult_125_G4_A_not_8_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_8_0_port);
   mult_125_G4_AN2_7_15 : nor2 port map( a => mult_125_G4_A_notx_7_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_7_15_port);
   mult_125_G4_AN1_7_14 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_7_14_port);
   mult_125_G4_AN1_7_13 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_7_13_port);
   mult_125_G4_AN1_7_12 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_7_12_port);
   mult_125_G4_AN1_7_11 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_7_11_port);
   mult_125_G4_AN1_7_10 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_7_10_port);
   mult_125_G4_AN1_7_9 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_7_9_port);
   mult_125_G4_AN1_7_8 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_7_8_port);
   mult_125_G4_AN1_7_7 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_7_7_port);
   mult_125_G4_AN1_7_6 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_7_6_port);
   mult_125_G4_AN1_7_5 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_7_5_port);
   mult_125_G4_AN1_7_4 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_7_4_port);
   mult_125_G4_AN1_7_3 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_7_3_port);
   mult_125_G4_AN1_7_2 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_7_2_port);
   mult_125_G4_AN1_7_1 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_7_1_port);
   mult_125_G4_AN1_7_0_0 : nor2 port map( a => mult_125_G4_A_not_7_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_7_0_port);
   mult_125_G4_AN2_6_15 : nor2 port map( a => mult_125_G4_A_notx_6_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_6_15_port);
   mult_125_G4_AN1_6_14 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_6_14_port);
   mult_125_G4_AN1_6_13 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_6_13_port);
   mult_125_G4_AN1_6_12 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_6_12_port);
   mult_125_G4_AN1_6_11 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_6_11_port);
   mult_125_G4_AN1_6_10 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_6_10_port);
   mult_125_G4_AN1_6_9 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_6_9_port);
   mult_125_G4_AN1_6_8 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_6_8_port);
   mult_125_G4_AN1_6_7 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_6_7_port);
   mult_125_G4_AN1_6_6 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_6_6_port);
   mult_125_G4_AN1_6_5 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_6_5_port);
   mult_125_G4_AN1_6_4 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_6_4_port);
   mult_125_G4_AN1_6_3 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_6_3_port);
   mult_125_G4_AN1_6_2 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_6_2_port);
   mult_125_G4_AN1_6_1 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_6_1_port);
   mult_125_G4_AN1_6_0_0 : nor2 port map( a => mult_125_G4_A_not_6_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_6_0_port);
   mult_125_G4_AN2_5_15 : nor2 port map( a => mult_125_G4_A_notx_5_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_5_15_port);
   mult_125_G4_AN1_5_14 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_5_14_port);
   mult_125_G4_AN1_5_13 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_5_13_port);
   mult_125_G4_AN1_5_12 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_5_12_port);
   mult_125_G4_AN1_5_11 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_5_11_port);
   mult_125_G4_AN1_5_10 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_5_10_port);
   mult_125_G4_AN1_5_9 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_5_9_port);
   mult_125_G4_AN1_5_8 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_5_8_port);
   mult_125_G4_AN1_5_7 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_5_7_port);
   mult_125_G4_AN1_5_6 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_5_6_port);
   mult_125_G4_AN1_5_5 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_5_5_port);
   mult_125_G4_AN1_5_4 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_5_4_port);
   mult_125_G4_AN1_5_3 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_5_3_port);
   mult_125_G4_AN1_5_2 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_5_2_port);
   mult_125_G4_AN1_5_1 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_5_1_port);
   mult_125_G4_AN1_5_0_0 : nor2 port map( a => mult_125_G4_A_not_5_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_5_0_port);
   mult_125_G4_AN2_4_15 : nor2 port map( a => mult_125_G4_A_notx_4_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_4_15_port);
   mult_125_G4_AN1_4_14 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_4_14_port);
   mult_125_G4_AN1_4_13 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_4_13_port);
   mult_125_G4_AN1_4_12 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_4_12_port);
   mult_125_G4_AN1_4_11 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_4_11_port);
   mult_125_G4_AN1_4_10 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_4_10_port);
   mult_125_G4_AN1_4_9 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_4_9_port);
   mult_125_G4_AN1_4_8 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_4_8_port);
   mult_125_G4_AN1_4_7 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_4_7_port);
   mult_125_G4_AN1_4_6 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_4_6_port);
   mult_125_G4_AN1_4_5 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_4_5_port);
   mult_125_G4_AN1_4_4 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_4_4_port);
   mult_125_G4_AN1_4_3 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_4_3_port);
   mult_125_G4_AN1_4_2 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_4_2_port);
   mult_125_G4_AN1_4_1 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_4_1_port);
   mult_125_G4_AN1_4_0_0 : nor2 port map( a => mult_125_G4_A_not_4_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_4_0_port);
   mult_125_G4_AN2_3_15 : nor2 port map( a => mult_125_G4_A_notx_3_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_3_15_port);
   mult_125_G4_AN1_3_14 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_3_14_port);
   mult_125_G4_AN1_3_13 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_3_13_port);
   mult_125_G4_AN1_3_12 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_3_12_port);
   mult_125_G4_AN1_3_11 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_3_11_port);
   mult_125_G4_AN1_3_10 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_3_10_port);
   mult_125_G4_AN1_3_9 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_3_9_port);
   mult_125_G4_AN1_3_8 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_3_8_port);
   mult_125_G4_AN1_3_7 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_3_7_port);
   mult_125_G4_AN1_3_6 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_3_6_port);
   mult_125_G4_AN1_3_5 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_3_5_port);
   mult_125_G4_AN1_3_4 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_3_4_port);
   mult_125_G4_AN1_3_3 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_3_3_port);
   mult_125_G4_AN1_3_2 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_3_2_port);
   mult_125_G4_AN1_3_1 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_3_1_port);
   mult_125_G4_AN1_3_0_0 : nor2 port map( a => mult_125_G4_A_not_3_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_3_0_port);
   mult_125_G4_AN2_2_15 : nor2 port map( a => mult_125_G4_A_notx_2_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_2_15_port);
   mult_125_G4_AN1_2_14 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_2_14_port);
   mult_125_G4_AN1_2_13 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_2_13_port);
   mult_125_G4_AN1_2_12 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_2_12_port);
   mult_125_G4_AN1_2_11 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_2_11_port);
   mult_125_G4_AN1_2_10 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_2_10_port);
   mult_125_G4_AN1_2_9 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_2_9_port);
   mult_125_G4_AN1_2_8 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_2_8_port);
   mult_125_G4_AN1_2_7 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_2_7_port);
   mult_125_G4_AN1_2_6 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_2_6_port);
   mult_125_G4_AN1_2_5 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_2_5_port);
   mult_125_G4_AN1_2_4 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_2_4_port);
   mult_125_G4_AN1_2_3 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_2_3_port);
   mult_125_G4_AN1_2_2 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_2_2_port);
   mult_125_G4_AN1_2_1 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_2_1_port);
   mult_125_G4_AN1_2_0_0 : nor2 port map( a => mult_125_G4_A_not_2_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_2_0_port);
   mult_125_G4_AN2_1_15 : nor2 port map( a => mult_125_G4_A_notx_1_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_1_15_port);
   mult_125_G4_AN1_1_14 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_1_14_port);
   mult_125_G4_AN1_1_13 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_1_13_port);
   mult_125_G4_AN1_1_12 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_1_12_port);
   mult_125_G4_AN1_1_11 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_1_11_port);
   mult_125_G4_AN1_1_10 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_1_10_port);
   mult_125_G4_AN1_1_9 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_1_9_port);
   mult_125_G4_AN1_1_8 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_1_8_port);
   mult_125_G4_AN1_1_7 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_1_7_port);
   mult_125_G4_AN1_1_6 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_1_6_port);
   mult_125_G4_AN1_1_5 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_1_5_port);
   mult_125_G4_AN1_1_4 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_1_4_port);
   mult_125_G4_AN1_1_3 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_1_3_port);
   mult_125_G4_AN1_1_2 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_1_2_port);
   mult_125_G4_AN1_1_1 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_1_1_port);
   mult_125_G4_AN1_1_0_0 : nor2 port map( a => mult_125_G4_A_not_1_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_ab_1_0_port);
   mult_125_G4_AN2_0_15 : nor2 port map( a => mult_125_G4_A_notx_0_port, b => 
                           mult_125_G4_B_not_15_port, outb => 
                           mult_125_G4_ab_0_15_port);
   mult_125_G4_AN1_0_14 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_ab_0_14_port);
   mult_125_G4_AN1_0_13 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_ab_0_13_port);
   mult_125_G4_AN1_0_12 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_ab_0_12_port);
   mult_125_G4_AN1_0_11 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_ab_0_11_port);
   mult_125_G4_AN1_0_10 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_ab_0_10_port);
   mult_125_G4_AN1_0_9 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_ab_0_9_port);
   mult_125_G4_AN1_0_8 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_ab_0_8_port);
   mult_125_G4_AN1_0_7 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_ab_0_7_port);
   mult_125_G4_AN1_0_6 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_ab_0_6_port);
   mult_125_G4_AN1_0_5 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_ab_0_5_port);
   mult_125_G4_AN1_0_4 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_ab_0_4_port);
   mult_125_G4_AN1_0_3 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_ab_0_3_port);
   mult_125_G4_AN1_0_2 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_ab_0_2_port);
   mult_125_G4_AN1_0_1 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_ab_0_1_port);
   mult_125_G4_AN1_0_0_0 : nor2 port map( a => mult_125_G4_A_not_0_port, b => 
                           mult_125_G4_B_not_0_port, outb => 
                           multiplier_sigs_3_0_port);
   U267 : inv port map( inb => input_sample_mem_15_port, outb => n5911);
   U268 : inv port map( inb => coefficient_mem_array_2_15_port, outb => n5912);
   U269 : inv port map( inb => mult_125_G3_B_not_15_port, outb => n5913);
   U270 : inv port map( inb => mult_125_G3_A_not_15_port, outb => n5914);
   U271 : inv port map( inb => mult_125_G3_A_not_0_port, outb => 
                           mult_125_G3_A_notx_0_port);
   U272 : inv port map( inb => mult_125_G3_A_not_1_port, outb => 
                           mult_125_G3_A_notx_1_port);
   U273 : inv port map( inb => mult_125_G3_A_not_2_port, outb => 
                           mult_125_G3_A_notx_2_port);
   U274 : inv port map( inb => mult_125_G3_A_not_3_port, outb => 
                           mult_125_G3_A_notx_3_port);
   U275 : inv port map( inb => mult_125_G3_A_not_4_port, outb => 
                           mult_125_G3_A_notx_4_port);
   U276 : inv port map( inb => mult_125_G3_A_not_5_port, outb => 
                           mult_125_G3_A_notx_5_port);
   U277 : inv port map( inb => mult_125_G3_A_not_6_port, outb => 
                           mult_125_G3_A_notx_6_port);
   U278 : inv port map( inb => mult_125_G3_A_not_7_port, outb => 
                           mult_125_G3_A_notx_7_port);
   U279 : inv port map( inb => mult_125_G3_A_not_8_port, outb => 
                           mult_125_G3_A_notx_8_port);
   U280 : inv port map( inb => mult_125_G3_A_not_9_port, outb => 
                           mult_125_G3_A_notx_9_port);
   U281 : inv port map( inb => mult_125_G3_A_not_10_port, outb => 
                           mult_125_G3_A_notx_10_port);
   U282 : inv port map( inb => mult_125_G3_A_not_11_port, outb => 
                           mult_125_G3_A_notx_11_port);
   U283 : inv port map( inb => mult_125_G3_A_not_12_port, outb => 
                           mult_125_G3_A_notx_12_port);
   U284 : inv port map( inb => mult_125_G3_A_not_13_port, outb => 
                           mult_125_G3_A_notx_13_port);
   U285 : inv port map( inb => mult_125_G3_A_not_14_port, outb => 
                           mult_125_G3_A_notx_14_port);
   U286 : inv port map( inb => mult_125_G3_B_not_0_port, outb => 
                           mult_125_G3_B_notx_0_port);
   U287 : inv port map( inb => mult_125_G3_B_not_1_port, outb => 
                           mult_125_G3_B_notx_1_port);
   U288 : inv port map( inb => mult_125_G3_B_not_2_port, outb => 
                           mult_125_G3_B_notx_2_port);
   U289 : inv port map( inb => mult_125_G3_B_not_3_port, outb => 
                           mult_125_G3_B_notx_3_port);
   U290 : inv port map( inb => mult_125_G3_B_not_4_port, outb => 
                           mult_125_G3_B_notx_4_port);
   U291 : inv port map( inb => mult_125_G3_B_not_5_port, outb => 
                           mult_125_G3_B_notx_5_port);
   U292 : inv port map( inb => mult_125_G3_B_not_6_port, outb => 
                           mult_125_G3_B_notx_6_port);
   U293 : inv port map( inb => mult_125_G3_B_not_7_port, outb => 
                           mult_125_G3_B_notx_7_port);
   U294 : inv port map( inb => mult_125_G3_B_not_8_port, outb => 
                           mult_125_G3_B_notx_8_port);
   U295 : inv port map( inb => mult_125_G3_B_not_9_port, outb => 
                           mult_125_G3_B_notx_9_port);
   U296 : inv port map( inb => mult_125_G3_B_not_10_port, outb => 
                           mult_125_G3_B_notx_10_port);
   U297 : inv port map( inb => mult_125_G3_B_not_11_port, outb => 
                           mult_125_G3_B_notx_11_port);
   U298 : inv port map( inb => mult_125_G3_B_not_12_port, outb => 
                           mult_125_G3_B_notx_12_port);
   U299 : inv port map( inb => mult_125_G3_B_not_13_port, outb => 
                           mult_125_G3_B_notx_13_port);
   U300 : inv port map( inb => mult_125_G3_B_not_14_port, outb => 
                           mult_125_G3_B_notx_14_port);
   U301 : inv port map( inb => input_sample_mem_15_port, outb => n5786);
   U302 : inv port map( inb => coefficient_mem_array_1_15_port, outb => n5787);
   U303 : inv port map( inb => mult_125_G2_B_not_15_port, outb => n5788);
   U304 : inv port map( inb => mult_125_G2_A_not_15_port, outb => n5789);
   U305 : inv port map( inb => mult_125_G2_A_not_0_port, outb => 
                           mult_125_G2_A_notx_0_port);
   U306 : inv port map( inb => mult_125_G2_A_not_1_port, outb => 
                           mult_125_G2_A_notx_1_port);
   U307 : inv port map( inb => mult_125_G2_A_not_2_port, outb => 
                           mult_125_G2_A_notx_2_port);
   U308 : inv port map( inb => mult_125_G2_A_not_3_port, outb => 
                           mult_125_G2_A_notx_3_port);
   U309 : inv port map( inb => mult_125_G2_A_not_4_port, outb => 
                           mult_125_G2_A_notx_4_port);
   U310 : inv port map( inb => mult_125_G2_A_not_5_port, outb => 
                           mult_125_G2_A_notx_5_port);
   U311 : inv port map( inb => mult_125_G2_A_not_6_port, outb => 
                           mult_125_G2_A_notx_6_port);
   U312 : inv port map( inb => mult_125_G2_A_not_7_port, outb => 
                           mult_125_G2_A_notx_7_port);
   U313 : inv port map( inb => mult_125_G2_A_not_8_port, outb => 
                           mult_125_G2_A_notx_8_port);
   U314 : inv port map( inb => mult_125_G2_A_not_9_port, outb => 
                           mult_125_G2_A_notx_9_port);
   U315 : inv port map( inb => mult_125_G2_A_not_10_port, outb => 
                           mult_125_G2_A_notx_10_port);
   U316 : inv port map( inb => mult_125_G2_A_not_11_port, outb => 
                           mult_125_G2_A_notx_11_port);
   U317 : inv port map( inb => mult_125_G2_A_not_12_port, outb => 
                           mult_125_G2_A_notx_12_port);
   U318 : inv port map( inb => mult_125_G2_A_not_13_port, outb => 
                           mult_125_G2_A_notx_13_port);
   U319 : inv port map( inb => mult_125_G2_A_not_14_port, outb => 
                           mult_125_G2_A_notx_14_port);
   U320 : inv port map( inb => mult_125_G2_B_not_0_port, outb => 
                           mult_125_G2_B_notx_0_port);
   U321 : inv port map( inb => mult_125_G2_B_not_1_port, outb => 
                           mult_125_G2_B_notx_1_port);
   U322 : inv port map( inb => mult_125_G2_B_not_2_port, outb => 
                           mult_125_G2_B_notx_2_port);
   U323 : inv port map( inb => mult_125_G2_B_not_3_port, outb => 
                           mult_125_G2_B_notx_3_port);
   U324 : inv port map( inb => mult_125_G2_B_not_4_port, outb => 
                           mult_125_G2_B_notx_4_port);
   U325 : inv port map( inb => mult_125_G2_B_not_5_port, outb => 
                           mult_125_G2_B_notx_5_port);
   U326 : inv port map( inb => mult_125_G2_B_not_6_port, outb => 
                           mult_125_G2_B_notx_6_port);
   U327 : inv port map( inb => mult_125_G2_B_not_7_port, outb => 
                           mult_125_G2_B_notx_7_port);
   U328 : inv port map( inb => mult_125_G2_B_not_8_port, outb => 
                           mult_125_G2_B_notx_8_port);
   U329 : inv port map( inb => mult_125_G2_B_not_9_port, outb => 
                           mult_125_G2_B_notx_9_port);
   U330 : inv port map( inb => mult_125_G2_B_not_10_port, outb => 
                           mult_125_G2_B_notx_10_port);
   U331 : inv port map( inb => mult_125_G2_B_not_11_port, outb => 
                           mult_125_G2_B_notx_11_port);
   U332 : inv port map( inb => mult_125_G2_B_not_12_port, outb => 
                           mult_125_G2_B_notx_12_port);
   U333 : inv port map( inb => mult_125_G2_B_not_13_port, outb => 
                           mult_125_G2_B_notx_13_port);
   U334 : inv port map( inb => mult_125_G2_B_not_14_port, outb => 
                           mult_125_G2_B_notx_14_port);
   U335 : inv port map( inb => input_sample_mem_15_port, outb => n5661);
   U336 : inv port map( inb => coefficient_mem_array_0_15_port, outb => n5662);
   U337 : inv port map( inb => mult_125_B_not_15_port, outb => n5663);
   U338 : inv port map( inb => mult_125_A_not_15_port, outb => n5664);
   U339 : inv port map( inb => mult_125_A_not_0_port, outb => 
                           mult_125_A_notx_0_port);
   U340 : inv port map( inb => mult_125_A_not_1_port, outb => 
                           mult_125_A_notx_1_port);
   U341 : inv port map( inb => mult_125_A_not_2_port, outb => 
                           mult_125_A_notx_2_port);
   U342 : inv port map( inb => mult_125_A_not_3_port, outb => 
                           mult_125_A_notx_3_port);
   U343 : inv port map( inb => mult_125_A_not_4_port, outb => 
                           mult_125_A_notx_4_port);
   U344 : inv port map( inb => mult_125_A_not_5_port, outb => 
                           mult_125_A_notx_5_port);
   U345 : inv port map( inb => mult_125_A_not_6_port, outb => 
                           mult_125_A_notx_6_port);
   U346 : inv port map( inb => mult_125_A_not_7_port, outb => 
                           mult_125_A_notx_7_port);
   U347 : inv port map( inb => mult_125_A_not_8_port, outb => 
                           mult_125_A_notx_8_port);
   U348 : inv port map( inb => mult_125_A_not_9_port, outb => 
                           mult_125_A_notx_9_port);
   U349 : inv port map( inb => mult_125_A_not_10_port, outb => 
                           mult_125_A_notx_10_port);
   U350 : inv port map( inb => mult_125_A_not_11_port, outb => 
                           mult_125_A_notx_11_port);
   U351 : inv port map( inb => mult_125_A_not_12_port, outb => 
                           mult_125_A_notx_12_port);
   U352 : inv port map( inb => mult_125_A_not_13_port, outb => 
                           mult_125_A_notx_13_port);
   U353 : inv port map( inb => mult_125_A_not_14_port, outb => 
                           mult_125_A_notx_14_port);
   U354 : inv port map( inb => mult_125_B_not_0_port, outb => 
                           mult_125_B_notx_0_port);
   U355 : inv port map( inb => mult_125_B_not_1_port, outb => 
                           mult_125_B_notx_1_port);
   U356 : inv port map( inb => mult_125_B_not_2_port, outb => 
                           mult_125_B_notx_2_port);
   U357 : inv port map( inb => mult_125_B_not_3_port, outb => 
                           mult_125_B_notx_3_port);
   U358 : inv port map( inb => mult_125_B_not_4_port, outb => 
                           mult_125_B_notx_4_port);
   U359 : inv port map( inb => mult_125_B_not_5_port, outb => 
                           mult_125_B_notx_5_port);
   U360 : inv port map( inb => mult_125_B_not_6_port, outb => 
                           mult_125_B_notx_6_port);
   U361 : inv port map( inb => mult_125_B_not_7_port, outb => 
                           mult_125_B_notx_7_port);
   U362 : inv port map( inb => mult_125_B_not_8_port, outb => 
                           mult_125_B_notx_8_port);
   U363 : inv port map( inb => mult_125_B_not_9_port, outb => 
                           mult_125_B_notx_9_port);
   U364 : inv port map( inb => mult_125_B_not_10_port, outb => 
                           mult_125_B_notx_10_port);
   U365 : inv port map( inb => mult_125_B_not_11_port, outb => 
                           mult_125_B_notx_11_port);
   U366 : inv port map( inb => mult_125_B_not_12_port, outb => 
                           mult_125_B_notx_12_port);
   U367 : inv port map( inb => mult_125_B_not_13_port, outb => 
                           mult_125_B_notx_13_port);
   U368 : inv port map( inb => mult_125_B_not_14_port, outb => 
                           mult_125_B_notx_14_port);
   U369 : inv port map( inb => input_sample_mem_15_port, outb => n5536);
   U370 : inv port map( inb => coefficient_mem_array_3_15_port, outb => n5537);
   U371 : inv port map( inb => mult_125_G4_B_not_15_port, outb => n5538);
   U372 : inv port map( inb => mult_125_G4_A_not_15_port, outb => n5539);
   U373 : inv port map( inb => mult_125_G4_A_not_0_port, outb => 
                           mult_125_G4_A_notx_0_port);
   U374 : inv port map( inb => mult_125_G4_A_not_1_port, outb => 
                           mult_125_G4_A_notx_1_port);
   U375 : inv port map( inb => mult_125_G4_A_not_2_port, outb => 
                           mult_125_G4_A_notx_2_port);
   U376 : inv port map( inb => mult_125_G4_A_not_3_port, outb => 
                           mult_125_G4_A_notx_3_port);
   U377 : inv port map( inb => mult_125_G4_A_not_4_port, outb => 
                           mult_125_G4_A_notx_4_port);
   U378 : inv port map( inb => mult_125_G4_A_not_5_port, outb => 
                           mult_125_G4_A_notx_5_port);
   U379 : inv port map( inb => mult_125_G4_A_not_6_port, outb => 
                           mult_125_G4_A_notx_6_port);
   U380 : inv port map( inb => mult_125_G4_A_not_7_port, outb => 
                           mult_125_G4_A_notx_7_port);
   U381 : inv port map( inb => mult_125_G4_A_not_8_port, outb => 
                           mult_125_G4_A_notx_8_port);
   U382 : inv port map( inb => mult_125_G4_A_not_9_port, outb => 
                           mult_125_G4_A_notx_9_port);
   U383 : inv port map( inb => mult_125_G4_A_not_10_port, outb => 
                           mult_125_G4_A_notx_10_port);
   U384 : inv port map( inb => mult_125_G4_A_not_11_port, outb => 
                           mult_125_G4_A_notx_11_port);
   U385 : inv port map( inb => mult_125_G4_A_not_12_port, outb => 
                           mult_125_G4_A_notx_12_port);
   U386 : inv port map( inb => mult_125_G4_A_not_13_port, outb => 
                           mult_125_G4_A_notx_13_port);
   U387 : inv port map( inb => mult_125_G4_A_not_14_port, outb => 
                           mult_125_G4_A_notx_14_port);
   U388 : inv port map( inb => mult_125_G4_B_not_0_port, outb => 
                           mult_125_G4_B_notx_0_port);
   U389 : inv port map( inb => mult_125_G4_B_not_1_port, outb => 
                           mult_125_G4_B_notx_1_port);
   U390 : inv port map( inb => mult_125_G4_B_not_2_port, outb => 
                           mult_125_G4_B_notx_2_port);
   U391 : inv port map( inb => mult_125_G4_B_not_3_port, outb => 
                           mult_125_G4_B_notx_3_port);
   U392 : inv port map( inb => mult_125_G4_B_not_4_port, outb => 
                           mult_125_G4_B_notx_4_port);
   U393 : inv port map( inb => mult_125_G4_B_not_5_port, outb => 
                           mult_125_G4_B_notx_5_port);
   U394 : inv port map( inb => mult_125_G4_B_not_6_port, outb => 
                           mult_125_G4_B_notx_6_port);
   U395 : inv port map( inb => mult_125_G4_B_not_7_port, outb => 
                           mult_125_G4_B_notx_7_port);
   U396 : inv port map( inb => mult_125_G4_B_not_8_port, outb => 
                           mult_125_G4_B_notx_8_port);
   U397 : inv port map( inb => mult_125_G4_B_not_9_port, outb => 
                           mult_125_G4_B_notx_9_port);
   U398 : inv port map( inb => mult_125_G4_B_not_10_port, outb => 
                           mult_125_G4_B_notx_10_port);
   U399 : inv port map( inb => mult_125_G4_B_not_11_port, outb => 
                           mult_125_G4_B_notx_11_port);
   U400 : inv port map( inb => mult_125_G4_B_not_12_port, outb => 
                           mult_125_G4_B_notx_12_port);
   U401 : inv port map( inb => mult_125_G4_B_not_13_port, outb => 
                           mult_125_G4_B_notx_13_port);
   U402 : inv port map( inb => mult_125_G4_B_not_14_port, outb => 
                           mult_125_G4_B_notx_14_port);
   U403 : inv port map( inb => n5540, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_0_0_port);
   U404 : inv port map( inb => n5660, outb => mult_125_G4_FS_1_C_1_4_0_port);
   U405 : inv port map( inb => n5665, outb => mult_125_FS_1_TEMP_P_0_0_0_port);
   U406 : inv port map( inb => n5785, outb => mult_125_FS_1_C_1_4_0_port);
   U407 : inv port map( inb => n5790, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_0_0_port);
   U408 : inv port map( inb => n5910, outb => mult_125_G2_FS_1_C_1_4_0_port);
   U409 : inv port map( inb => n5915, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_0_0_port);
   U410 : inv port map( inb => n6035, outb => mult_125_G3_FS_1_C_1_4_0_port);
   U411 : inv port map( inb => mult_125_FS_1_TEMP_P_0_0_0_port, outb => n5666);
   U412 : inv port map( inb => n5667, outb => mult_125_FS_1_P_0_0_1_port);
   U413 : inv port map( inb => mult_125_FS_1_P_0_0_1_port, outb => n5668);
   U414 : inv port map( inb => n5669, outb => mult_125_FS_1_P_0_0_2_port);
   U415 : inv port map( inb => mult_125_FS_1_P_0_0_2_port, outb => n5670);
   U416 : inv port map( inb => n5671, outb => mult_125_FS_1_P_0_0_3_port);
   U417 : inv port map( inb => mult_125_FS_1_P_0_0_3_port, outb => n5672);
   U418 : inv port map( inb => n5673, outb => mult_125_FS_1_TEMP_P_0_1_0_port);
   U419 : inv port map( inb => mult_125_FS_1_TEMP_P_0_1_0_port, outb => n5674);
   U420 : inv port map( inb => n5675, outb => mult_125_FS_1_P_0_1_1_port);
   U421 : inv port map( inb => mult_125_FS_1_P_0_1_1_port, outb => n5676);
   U422 : inv port map( inb => n5677, outb => mult_125_FS_1_P_0_1_2_port);
   U423 : inv port map( inb => mult_125_FS_1_P_0_1_2_port, outb => n5678);
   U424 : inv port map( inb => n5679, outb => mult_125_FS_1_P_0_1_3_port);
   U425 : inv port map( inb => mult_125_FS_1_P_0_1_3_port, outb => n5680);
   U426 : inv port map( inb => n5681, outb => mult_125_FS_1_TEMP_P_0_2_0_port);
   U427 : inv port map( inb => mult_125_FS_1_TEMP_P_0_2_0_port, outb => n5682);
   U428 : inv port map( inb => n5683, outb => mult_125_FS_1_P_0_2_1_port);
   U429 : inv port map( inb => mult_125_FS_1_P_0_2_1_port, outb => n5684);
   U430 : inv port map( inb => n5685, outb => mult_125_FS_1_P_0_2_2_port);
   U431 : inv port map( inb => mult_125_FS_1_P_0_2_2_port, outb => n5686);
   U432 : inv port map( inb => n5687, outb => mult_125_FS_1_P_0_2_3_port);
   U433 : inv port map( inb => mult_125_FS_1_P_0_2_3_port, outb => n5688);
   U434 : inv port map( inb => n5775, outb => mult_125_FS_1_G_2_0_0_port);
   U435 : inv port map( inb => n5689, outb => mult_125_FS_1_TEMP_P_0_3_0_port);
   U436 : inv port map( inb => mult_125_FS_1_TEMP_P_0_3_0_port, outb => n5690);
   U437 : inv port map( inb => n5691, outb => mult_125_FS_1_P_0_3_1_port);
   U438 : inv port map( inb => mult_125_FS_1_P_0_3_1_port, outb => n5692);
   U439 : inv port map( inb => mult_125_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_FS_1_C_1_3_3_port);
   U440 : inv port map( inb => mult_125_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_FS_1_TEMP_G_0_3_2_port);
   U441 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_0_0_port, outb => 
                           n5791);
   U442 : inv port map( inb => n5792, outb => mult_125_G2_FS_1_P_0_0_1_port);
   U443 : inv port map( inb => mult_125_G2_FS_1_P_0_0_1_port, outb => n5793);
   U444 : inv port map( inb => n5794, outb => mult_125_G2_FS_1_P_0_0_2_port);
   U445 : inv port map( inb => mult_125_G2_FS_1_P_0_0_2_port, outb => n5795);
   U446 : inv port map( inb => n5796, outb => mult_125_G2_FS_1_P_0_0_3_port);
   U447 : inv port map( inb => mult_125_G2_FS_1_P_0_0_3_port, outb => n5797);
   U448 : inv port map( inb => n5798, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_1_0_port);
   U449 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_1_0_port, outb => 
                           n5799);
   U450 : inv port map( inb => n5800, outb => mult_125_G2_FS_1_P_0_1_1_port);
   U451 : inv port map( inb => mult_125_G2_FS_1_P_0_1_1_port, outb => n5801);
   U452 : inv port map( inb => n5802, outb => mult_125_G2_FS_1_P_0_1_2_port);
   U453 : inv port map( inb => mult_125_G2_FS_1_P_0_1_2_port, outb => n5803);
   U454 : inv port map( inb => n5804, outb => mult_125_G2_FS_1_P_0_1_3_port);
   U455 : inv port map( inb => mult_125_G2_FS_1_P_0_1_3_port, outb => n5805);
   U456 : inv port map( inb => n5806, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_2_0_port);
   U457 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_2_0_port, outb => 
                           n5807);
   U458 : inv port map( inb => n5808, outb => mult_125_G2_FS_1_P_0_2_1_port);
   U459 : inv port map( inb => mult_125_G2_FS_1_P_0_2_1_port, outb => n5809);
   U460 : inv port map( inb => n5810, outb => mult_125_G2_FS_1_P_0_2_2_port);
   U461 : inv port map( inb => mult_125_G2_FS_1_P_0_2_2_port, outb => n5811);
   U462 : inv port map( inb => n5812, outb => mult_125_G2_FS_1_P_0_2_3_port);
   U463 : inv port map( inb => mult_125_G2_FS_1_P_0_2_3_port, outb => n5813);
   U464 : inv port map( inb => n5900, outb => mult_125_G2_FS_1_G_2_0_0_port);
   U465 : inv port map( inb => n5814, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_3_0_port);
   U466 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_3_0_port, outb => 
                           n5815);
   U467 : inv port map( inb => n5816, outb => mult_125_G2_FS_1_P_0_3_1_port);
   U468 : inv port map( inb => mult_125_G2_FS_1_P_0_3_1_port, outb => n5817);
   U469 : inv port map( inb => mult_125_G2_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G2_FS_1_C_1_3_3_port);
   U470 : inv port map( inb => mult_125_G2_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G2_FS_1_TEMP_G_0_3_2_port);
   U471 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_0_0_port, outb => 
                           n5916);
   U472 : inv port map( inb => n5917, outb => mult_125_G3_FS_1_P_0_0_1_port);
   U473 : inv port map( inb => mult_125_G3_FS_1_P_0_0_1_port, outb => n5918);
   U474 : inv port map( inb => n5919, outb => mult_125_G3_FS_1_P_0_0_2_port);
   U475 : inv port map( inb => mult_125_G3_FS_1_P_0_0_2_port, outb => n5920);
   U476 : inv port map( inb => n5921, outb => mult_125_G3_FS_1_P_0_0_3_port);
   U477 : inv port map( inb => mult_125_G3_FS_1_P_0_0_3_port, outb => n5922);
   U478 : inv port map( inb => n5923, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_1_0_port);
   U479 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_1_0_port, outb => 
                           n5924);
   U480 : inv port map( inb => n5925, outb => mult_125_G3_FS_1_P_0_1_1_port);
   U481 : inv port map( inb => mult_125_G3_FS_1_P_0_1_1_port, outb => n5926);
   U482 : inv port map( inb => n5927, outb => mult_125_G3_FS_1_P_0_1_2_port);
   U483 : inv port map( inb => mult_125_G3_FS_1_P_0_1_2_port, outb => n5928);
   U484 : inv port map( inb => n5929, outb => mult_125_G3_FS_1_P_0_1_3_port);
   U485 : inv port map( inb => mult_125_G3_FS_1_P_0_1_3_port, outb => n5930);
   U486 : inv port map( inb => n5931, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_2_0_port);
   U487 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_2_0_port, outb => 
                           n5932);
   U488 : inv port map( inb => n5933, outb => mult_125_G3_FS_1_P_0_2_1_port);
   U489 : inv port map( inb => mult_125_G3_FS_1_P_0_2_1_port, outb => n5934);
   U490 : inv port map( inb => n5935, outb => mult_125_G3_FS_1_P_0_2_2_port);
   U491 : inv port map( inb => mult_125_G3_FS_1_P_0_2_2_port, outb => n5936);
   U492 : inv port map( inb => n5937, outb => mult_125_G3_FS_1_P_0_2_3_port);
   U493 : inv port map( inb => mult_125_G3_FS_1_P_0_2_3_port, outb => n5938);
   U494 : inv port map( inb => n6025, outb => mult_125_G3_FS_1_G_2_0_0_port);
   U495 : inv port map( inb => n5939, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_3_0_port);
   U496 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_3_0_port, outb => 
                           n5940);
   U497 : inv port map( inb => n5941, outb => mult_125_G3_FS_1_P_0_3_1_port);
   U498 : inv port map( inb => mult_125_G3_FS_1_P_0_3_1_port, outb => n5942);
   U499 : inv port map( inb => mult_125_G3_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G3_FS_1_C_1_3_3_port);
   U500 : inv port map( inb => mult_125_G3_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G3_FS_1_TEMP_G_0_3_2_port);
   U501 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_0_0_port, outb => 
                           n5541);
   U502 : inv port map( inb => n5542, outb => mult_125_G4_FS_1_P_0_0_1_port);
   U503 : inv port map( inb => mult_125_G4_FS_1_P_0_0_1_port, outb => n5543);
   U504 : inv port map( inb => n5544, outb => mult_125_G4_FS_1_P_0_0_2_port);
   U505 : inv port map( inb => mult_125_G4_FS_1_P_0_0_2_port, outb => n5545);
   U506 : inv port map( inb => n5546, outb => mult_125_G4_FS_1_P_0_0_3_port);
   U507 : inv port map( inb => mult_125_G4_FS_1_P_0_0_3_port, outb => n5547);
   U508 : inv port map( inb => n5548, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_1_0_port);
   U509 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_1_0_port, outb => 
                           n5549);
   U510 : inv port map( inb => n5550, outb => mult_125_G4_FS_1_P_0_1_1_port);
   U511 : inv port map( inb => mult_125_G4_FS_1_P_0_1_1_port, outb => n5551);
   U512 : inv port map( inb => n5552, outb => mult_125_G4_FS_1_P_0_1_2_port);
   U513 : inv port map( inb => mult_125_G4_FS_1_P_0_1_2_port, outb => n5553);
   U514 : inv port map( inb => n5554, outb => mult_125_G4_FS_1_P_0_1_3_port);
   U515 : inv port map( inb => mult_125_G4_FS_1_P_0_1_3_port, outb => n5555);
   U516 : inv port map( inb => n5556, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_2_0_port);
   U517 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_2_0_port, outb => 
                           n5557);
   U518 : inv port map( inb => n5558, outb => mult_125_G4_FS_1_P_0_2_1_port);
   U519 : inv port map( inb => mult_125_G4_FS_1_P_0_2_1_port, outb => n5559);
   U520 : inv port map( inb => n5560, outb => mult_125_G4_FS_1_P_0_2_2_port);
   U521 : inv port map( inb => mult_125_G4_FS_1_P_0_2_2_port, outb => n5561);
   U522 : inv port map( inb => n5562, outb => mult_125_G4_FS_1_P_0_2_3_port);
   U523 : inv port map( inb => mult_125_G4_FS_1_P_0_2_3_port, outb => n5563);
   U524 : inv port map( inb => n5650, outb => mult_125_G4_FS_1_G_2_0_0_port);
   U525 : inv port map( inb => n5564, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_3_0_port);
   U526 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_3_0_port, outb => 
                           n5565);
   U527 : inv port map( inb => n5566, outb => mult_125_G4_FS_1_P_0_3_1_port);
   U528 : inv port map( inb => mult_125_G4_FS_1_P_0_3_1_port, outb => n5567);
   U529 : inv port map( inb => mult_125_G4_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G4_FS_1_C_1_3_3_port);
   U530 : inv port map( inb => mult_125_G4_FS_1_G_n_int_0_3_2_port, outb => 
                           mult_125_G4_FS_1_TEMP_G_0_3_2_port);
   U531 : oai22 port map( a => mult_125_G4_QB, b => mult_125_G4_ab_15_15_port, 
                           c => mult_125_G4_QA, d => n240, outb => 
                           mult_125_G4_A1_29_port);
   U532 : nor2 port map( a => n241, b => n242, outb => mult_125_G4_A2_29_port);
   U533 : nor2 port map( a => n243, b => n244, outb => mult_125_G4_A2_28_port);
   U534 : nor2 port map( a => n245, b => n246, outb => mult_125_G4_A2_27_port);
   U535 : nor2 port map( a => n247, b => n248, outb => mult_125_G4_A2_26_port);
   U536 : nor2 port map( a => n249, b => n250, outb => mult_125_G4_A2_25_port);
   U537 : nor2 port map( a => n251, b => n252, outb => mult_125_G4_A2_24_port);
   U538 : nor2 port map( a => n253, b => n254, outb => mult_125_G4_A2_23_port);
   U539 : nor2 port map( a => n255, b => n256, outb => mult_125_G4_A2_22_port);
   U540 : nor2 port map( a => n257, b => n258, outb => mult_125_G4_A2_21_port);
   U541 : nor2 port map( a => n259, b => n260, outb => mult_125_G4_A2_20_port);
   U542 : nor2 port map( a => n261, b => n262, outb => mult_125_G4_A2_19_port);
   U543 : nor2 port map( a => n263, b => n264, outb => mult_125_G4_A2_18_port);
   U544 : nand2 port map( a => n266, b => n267, outb => n265);
   U545 : nor2 port map( a => n268, b => n269, outb => mult_125_G4_A2_16_port);
   U546 : nor2 port map( a => n270, b => n271, outb => mult_125_G4_A2_15_port);
   U547 : oai22 port map( a => n272, b => n273, c => n274, d => n275, outb => 
                           mult_125_G4_A2_14_port);
   U548 : oai22 port map( a => mult_125_QB, b => mult_125_ab_15_15_port, c => 
                           mult_125_QA, d => n276, outb => mult_125_A1_29_port)
                           ;
   U549 : nor2 port map( a => n277, b => n278, outb => mult_125_A2_29_port);
   U550 : nor2 port map( a => n279, b => n280, outb => mult_125_A2_28_port);
   U551 : nor2 port map( a => n281, b => n282, outb => mult_125_A2_27_port);
   U552 : nor2 port map( a => n283, b => n284, outb => mult_125_A2_26_port);
   U553 : nor2 port map( a => n285, b => n286, outb => mult_125_A2_25_port);
   U554 : nor2 port map( a => n287, b => n288, outb => mult_125_A2_24_port);
   U555 : nor2 port map( a => n289, b => n290, outb => mult_125_A2_23_port);
   U556 : nor2 port map( a => n291, b => n292, outb => mult_125_A2_22_port);
   U557 : nor2 port map( a => n293, b => n294, outb => mult_125_A2_21_port);
   U558 : nor2 port map( a => n295, b => n296, outb => mult_125_A2_20_port);
   U559 : nor2 port map( a => n297, b => n298, outb => mult_125_A2_19_port);
   U560 : nor2 port map( a => n299, b => n300, outb => mult_125_A2_18_port);
   U561 : nand2 port map( a => n302, b => n303, outb => n301);
   U562 : nor2 port map( a => n304, b => n305, outb => mult_125_A2_16_port);
   U563 : nor2 port map( a => n306, b => n307, outb => mult_125_A2_15_port);
   U564 : oai22 port map( a => n308, b => n309, c => n310, d => n311, outb => 
                           mult_125_A2_14_port);
   U565 : oai22 port map( a => mult_125_G2_QB, b => mult_125_G2_ab_15_15_port, 
                           c => mult_125_G2_QA, d => n312, outb => 
                           mult_125_G2_A1_29_port);
   U566 : nor2 port map( a => n313, b => n314, outb => mult_125_G2_A2_29_port);
   U567 : nor2 port map( a => n315, b => n316, outb => mult_125_G2_A2_28_port);
   U568 : nor2 port map( a => n317, b => n318, outb => mult_125_G2_A2_27_port);
   U569 : nor2 port map( a => n319, b => n320, outb => mult_125_G2_A2_26_port);
   U570 : nor2 port map( a => n321, b => n322, outb => mult_125_G2_A2_25_port);
   U571 : nor2 port map( a => n323, b => n324, outb => mult_125_G2_A2_24_port);
   U572 : nor2 port map( a => n325, b => n326, outb => mult_125_G2_A2_23_port);
   U573 : nor2 port map( a => n327, b => n328, outb => mult_125_G2_A2_22_port);
   U574 : nor2 port map( a => n329, b => n330, outb => mult_125_G2_A2_21_port);
   U575 : nor2 port map( a => n331, b => n332, outb => mult_125_G2_A2_20_port);
   U576 : nor2 port map( a => n333, b => n334, outb => mult_125_G2_A2_19_port);
   U577 : nor2 port map( a => n335, b => n336, outb => mult_125_G2_A2_18_port);
   U578 : nand2 port map( a => n338, b => n339, outb => n337);
   U579 : nor2 port map( a => n340, b => n341, outb => mult_125_G2_A2_16_port);
   U580 : nor2 port map( a => n342, b => n343, outb => mult_125_G2_A2_15_port);
   U581 : oai22 port map( a => n344, b => n345, c => n346, d => n347, outb => 
                           mult_125_G2_A2_14_port);
   U582 : oai22 port map( a => mult_125_G3_QB, b => mult_125_G3_ab_15_15_port, 
                           c => mult_125_G3_QA, d => n348, outb => 
                           mult_125_G3_A1_29_port);
   U583 : nor2 port map( a => n349, b => n350, outb => mult_125_G3_A2_29_port);
   U584 : nor2 port map( a => n351, b => n352, outb => mult_125_G3_A2_28_port);
   U585 : nor2 port map( a => n353, b => n354, outb => mult_125_G3_A2_27_port);
   U586 : nor2 port map( a => n355, b => n356, outb => mult_125_G3_A2_26_port);
   U587 : nor2 port map( a => n357, b => n358, outb => mult_125_G3_A2_25_port);
   U588 : nor2 port map( a => n359, b => n360, outb => mult_125_G3_A2_24_port);
   U589 : nor2 port map( a => n361, b => n362, outb => mult_125_G3_A2_23_port);
   U590 : nor2 port map( a => n363, b => n364, outb => mult_125_G3_A2_22_port);
   U591 : nor2 port map( a => n365, b => n366, outb => mult_125_G3_A2_21_port);
   U592 : nor2 port map( a => n367, b => n368, outb => mult_125_G3_A2_20_port);
   U593 : nor2 port map( a => n369, b => n370, outb => mult_125_G3_A2_19_port);
   U594 : nor2 port map( a => n371, b => n372, outb => mult_125_G3_A2_18_port);
   U595 : nand2 port map( a => n374, b => n375, outb => n373);
   U596 : nor2 port map( a => n376, b => n377, outb => mult_125_G3_A2_16_port);
   U597 : nor2 port map( a => n378, b => n379, outb => mult_125_G3_A2_15_port);
   U598 : oai22 port map( a => n380, b => n381, c => n382, d => n383, outb => 
                           mult_125_G3_A2_14_port);
   U599 : nor2 port map( a => mult_125_G4_ab_1_15_port, b => 
                           mult_125_G4_ab_2_14_port, outb => n384);
   U600 : nor2 port map( a => mult_125_G4_ab_2_15_port, b => 
                           mult_125_G4_ab_3_14_port, outb => n385);
   U601 : nor2 port map( a => mult_125_G4_ab_3_15_port, b => 
                           mult_125_G4_ab_4_14_port, outb => n386);
   U602 : nor2 port map( a => mult_125_G4_ab_4_15_port, b => 
                           mult_125_G4_ab_5_14_port, outb => n387);
   U603 : nor2 port map( a => mult_125_G4_ab_5_15_port, b => 
                           mult_125_G4_ab_6_14_port, outb => n388);
   U604 : nor2 port map( a => mult_125_G4_ab_6_15_port, b => 
                           mult_125_G4_ab_7_14_port, outb => n389);
   U605 : nor2 port map( a => mult_125_G4_ab_7_15_port, b => 
                           mult_125_G4_ab_8_14_port, outb => n390);
   U606 : nor2 port map( a => mult_125_G4_ab_8_15_port, b => 
                           mult_125_G4_ab_9_14_port, outb => n391);
   U607 : nor2 port map( a => mult_125_G4_ab_9_15_port, b => 
                           mult_125_G4_ab_10_14_port, outb => n392);
   U608 : nor2 port map( a => mult_125_G4_ab_10_15_port, b => 
                           mult_125_G4_ab_11_14_port, outb => n393);
   U609 : nor2 port map( a => mult_125_G4_ab_11_15_port, b => 
                           mult_125_G4_ab_12_14_port, outb => n394);
   U610 : nor2 port map( a => mult_125_G4_ab_12_15_port, b => 
                           mult_125_G4_ab_13_14_port, outb => n395);
   U611 : nor2 port map( a => mult_125_G4_ab_13_15_port, b => 
                           mult_125_G4_ab_14_14_port, outb => n396);
   U612 : nor2 port map( a => mult_125_G4_ab_14_15_port, b => 
                           mult_125_G4_ab_15_14_port, outb => n397);
   U613 : nand2 port map( a => n399, b => n400, outb => n398);
   U614 : nand2 port map( a => n402, b => n403, outb => n401);
   U615 : nor2 port map( a => mult_125_G4_ab_4_13_port, b => n405, outb => n404
                           );
   U616 : nor2 port map( a => mult_125_G4_ab_5_13_port, b => n407, outb => n406
                           );
   U617 : nor2 port map( a => mult_125_G4_ab_6_13_port, b => n409, outb => n408
                           );
   U618 : nor2 port map( a => mult_125_G4_ab_7_13_port, b => n411, outb => n410
                           );
   U619 : nor2 port map( a => mult_125_G4_ab_8_13_port, b => n413, outb => n412
                           );
   U620 : nor2 port map( a => mult_125_G4_ab_9_13_port, b => n415, outb => n414
                           );
   U621 : nor2 port map( a => mult_125_G4_ab_10_13_port, b => n417, outb => 
                           n416);
   U622 : nor2 port map( a => mult_125_G4_ab_11_13_port, b => n419, outb => 
                           n418);
   U623 : nor2 port map( a => mult_125_G4_ab_12_13_port, b => n421, outb => 
                           n420);
   U624 : nor2 port map( a => mult_125_G4_ab_13_13_port, b => n423, outb => 
                           n422);
   U625 : nor2 port map( a => mult_125_G4_ab_14_13_port, b => n425, outb => 
                           n424);
   U626 : nor2 port map( a => mult_125_G4_ab_15_13_port, b => n427, outb => 
                           n426);
   U627 : nand2 port map( a => n429, b => n430, outb => n428);
   U628 : nor2 port map( a => mult_125_G4_ab_3_12_port, b => n432, outb => n431
                           );
   U629 : nor2 port map( a => mult_125_G4_ab_4_12_port, b => n434, outb => n433
                           );
   U630 : nor2 port map( a => mult_125_G4_ab_5_12_port, b => n436, outb => n435
                           );
   U631 : nor2 port map( a => mult_125_G4_ab_6_12_port, b => n438, outb => n437
                           );
   U632 : nor2 port map( a => mult_125_G4_ab_7_12_port, b => n440, outb => n439
                           );
   U633 : nor2 port map( a => mult_125_G4_ab_8_12_port, b => n442, outb => n441
                           );
   U634 : nor2 port map( a => mult_125_G4_ab_9_12_port, b => n444, outb => n443
                           );
   U635 : nor2 port map( a => mult_125_G4_ab_10_12_port, b => n446, outb => 
                           n445);
   U636 : nor2 port map( a => mult_125_G4_ab_11_12_port, b => n448, outb => 
                           n447);
   U637 : nor2 port map( a => mult_125_G4_ab_12_12_port, b => n450, outb => 
                           n449);
   U638 : nor2 port map( a => mult_125_G4_ab_13_12_port, b => n452, outb => 
                           n451);
   U639 : nor2 port map( a => mult_125_G4_ab_14_12_port, b => n454, outb => 
                           n453);
   U640 : nor2 port map( a => mult_125_G4_ab_15_12_port, b => n456, outb => 
                           n455);
   U641 : nand2 port map( a => n458, b => n459, outb => n457);
   U642 : nand2 port map( a => n461, b => n462, outb => n460);
   U643 : nor2 port map( a => mult_125_G4_ab_4_11_port, b => n464, outb => n463
                           );
   U644 : nor2 port map( a => mult_125_G4_ab_5_11_port, b => n466, outb => n465
                           );
   U645 : nor2 port map( a => mult_125_G4_ab_6_11_port, b => n468, outb => n467
                           );
   U646 : nor2 port map( a => mult_125_G4_ab_7_11_port, b => n470, outb => n469
                           );
   U647 : nor2 port map( a => mult_125_G4_ab_8_11_port, b => n472, outb => n471
                           );
   U648 : nor2 port map( a => mult_125_G4_ab_9_11_port, b => n474, outb => n473
                           );
   U649 : nor2 port map( a => mult_125_G4_ab_10_11_port, b => n476, outb => 
                           n475);
   U650 : nor2 port map( a => mult_125_G4_ab_11_11_port, b => n478, outb => 
                           n477);
   U651 : nor2 port map( a => mult_125_G4_ab_12_11_port, b => n480, outb => 
                           n479);
   U652 : nor2 port map( a => mult_125_G4_ab_13_11_port, b => n482, outb => 
                           n481);
   U653 : nor2 port map( a => mult_125_G4_ab_14_11_port, b => n484, outb => 
                           n483);
   U654 : nand2 port map( a => n486, b => n487, outb => n485);
   U655 : nand2 port map( a => n489, b => n490, outb => n488);
   U656 : nor2 port map( a => mult_125_G4_ab_3_10_port, b => n492, outb => n491
                           );
   U657 : nor2 port map( a => mult_125_G4_ab_4_10_port, b => n494, outb => n493
                           );
   U658 : nand2 port map( a => n496, b => n497, outb => n495);
   U659 : nor2 port map( a => mult_125_G4_ab_6_10_port, b => n499, outb => n498
                           );
   U660 : nor2 port map( a => mult_125_G4_ab_7_10_port, b => n501, outb => n500
                           );
   U661 : nor2 port map( a => mult_125_G4_ab_8_10_port, b => n503, outb => n502
                           );
   U662 : nor2 port map( a => mult_125_G4_ab_9_10_port, b => n505, outb => n504
                           );
   U663 : nor2 port map( a => mult_125_G4_ab_10_10_port, b => n507, outb => 
                           n506);
   U664 : nor2 port map( a => mult_125_G4_ab_11_10_port, b => n509, outb => 
                           n508);
   U665 : nor2 port map( a => mult_125_G4_ab_12_10_port, b => n511, outb => 
                           n510);
   U666 : nor2 port map( a => mult_125_G4_ab_13_10_port, b => n513, outb => 
                           n512);
   U667 : nor2 port map( a => mult_125_G4_ab_14_10_port, b => n515, outb => 
                           n514);
   U668 : nor2 port map( a => mult_125_G4_ab_15_10_port, b => n517, outb => 
                           n516);
   U669 : nand2 port map( a => n519, b => n520, outb => n518);
   U670 : nor2 port map( a => mult_125_G4_ab_3_9_port, b => n522, outb => n521)
                           ;
   U671 : nor2 port map( a => mult_125_G4_ab_4_9_port, b => n524, outb => n523)
                           ;
   U672 : nor2 port map( a => mult_125_G4_ab_5_9_port, b => n526, outb => n525)
                           ;
   U673 : nor2 port map( a => mult_125_G4_ab_6_9_port, b => n528, outb => n527)
                           ;
   U674 : nor2 port map( a => mult_125_G4_ab_7_9_port, b => n530, outb => n529)
                           ;
   U675 : nor2 port map( a => mult_125_G4_ab_8_9_port, b => n532, outb => n531)
                           ;
   U676 : nor2 port map( a => mult_125_G4_ab_9_9_port, b => n534, outb => n533)
                           ;
   U677 : nor2 port map( a => mult_125_G4_ab_10_9_port, b => n536, outb => n535
                           );
   U678 : nor2 port map( a => mult_125_G4_ab_11_9_port, b => n538, outb => n537
                           );
   U679 : nor2 port map( a => mult_125_G4_ab_12_9_port, b => n540, outb => n539
                           );
   U680 : nor2 port map( a => mult_125_G4_ab_13_9_port, b => n542, outb => n541
                           );
   U681 : nor2 port map( a => mult_125_G4_ab_14_9_port, b => n544, outb => n543
                           );
   U682 : nand2 port map( a => n546, b => n547, outb => n545);
   U683 : nand2 port map( a => n549, b => n550, outb => n548);
   U684 : nor2 port map( a => mult_125_G4_ab_3_8_port, b => n552, outb => n551)
                           ;
   U685 : nor2 port map( a => mult_125_G4_ab_4_8_port, b => n554, outb => n553)
                           ;
   U686 : nor2 port map( a => mult_125_G4_ab_5_8_port, b => n556, outb => n555)
                           ;
   U687 : nor2 port map( a => mult_125_G4_ab_6_8_port, b => n558, outb => n557)
                           ;
   U688 : nor2 port map( a => mult_125_G4_ab_7_8_port, b => n560, outb => n559)
                           ;
   U689 : nor2 port map( a => mult_125_G4_ab_8_8_port, b => n562, outb => n561)
                           ;
   U690 : nor2 port map( a => mult_125_G4_ab_9_8_port, b => n564, outb => n563)
                           ;
   U691 : nor2 port map( a => mult_125_G4_ab_10_8_port, b => n566, outb => n565
                           );
   U692 : nor2 port map( a => mult_125_G4_ab_11_8_port, b => n568, outb => n567
                           );
   U693 : nor2 port map( a => mult_125_G4_ab_12_8_port, b => n570, outb => n569
                           );
   U694 : nor2 port map( a => mult_125_G4_ab_13_8_port, b => n572, outb => n571
                           );
   U695 : nor2 port map( a => mult_125_G4_ab_14_8_port, b => n574, outb => n573
                           );
   U696 : nor2 port map( a => mult_125_G4_ab_15_8_port, b => n576, outb => n575
                           );
   U697 : nand2 port map( a => n578, b => n579, outb => n577);
   U698 : nand2 port map( a => n581, b => n582, outb => n580);
   U699 : nor2 port map( a => mult_125_G4_ab_4_7_port, b => n584, outb => n583)
                           ;
   U700 : nor2 port map( a => mult_125_G4_ab_5_7_port, b => n586, outb => n585)
                           ;
   U701 : nor2 port map( a => mult_125_G4_ab_6_7_port, b => n588, outb => n587)
                           ;
   U702 : nor2 port map( a => mult_125_G4_ab_7_7_port, b => n590, outb => n589)
                           ;
   U703 : nor2 port map( a => mult_125_G4_ab_8_7_port, b => n592, outb => n591)
                           ;
   U704 : nor2 port map( a => mult_125_G4_ab_9_7_port, b => n594, outb => n593)
                           ;
   U705 : nor2 port map( a => mult_125_G4_ab_10_7_port, b => n596, outb => n595
                           );
   U706 : nor2 port map( a => mult_125_G4_ab_11_7_port, b => n598, outb => n597
                           );
   U707 : nor2 port map( a => mult_125_G4_ab_12_7_port, b => n600, outb => n599
                           );
   U708 : nor2 port map( a => mult_125_G4_ab_13_7_port, b => n602, outb => n601
                           );
   U709 : nor2 port map( a => mult_125_G4_ab_14_7_port, b => n604, outb => n603
                           );
   U710 : nand2 port map( a => n606, b => n607, outb => n605);
   U711 : nand2 port map( a => n609, b => n610, outb => n608);
   U712 : nor2 port map( a => mult_125_G4_ab_3_6_port, b => n612, outb => n611)
                           ;
   U713 : nor2 port map( a => mult_125_G4_ab_4_6_port, b => n614, outb => n613)
                           ;
   U714 : nand2 port map( a => n616, b => n617, outb => n615);
   U715 : nor2 port map( a => mult_125_G4_ab_6_6_port, b => n619, outb => n618)
                           ;
   U716 : nor2 port map( a => mult_125_G4_ab_7_6_port, b => n621, outb => n620)
                           ;
   U717 : nor2 port map( a => mult_125_G4_ab_8_6_port, b => n623, outb => n622)
                           ;
   U718 : nand2 port map( a => n625, b => n626, outb => n624);
   U719 : nor2 port map( a => mult_125_G4_ab_10_6_port, b => n628, outb => n627
                           );
   U720 : nor2 port map( a => mult_125_G4_ab_11_6_port, b => n630, outb => n629
                           );
   U721 : nor2 port map( a => mult_125_G4_ab_12_6_port, b => n632, outb => n631
                           );
   U722 : nor2 port map( a => mult_125_G4_ab_13_6_port, b => n634, outb => n633
                           );
   U723 : nor2 port map( a => mult_125_G4_ab_14_6_port, b => n636, outb => n635
                           );
   U724 : nor2 port map( a => mult_125_G4_ab_15_6_port, b => n638, outb => n637
                           );
   U725 : nand2 port map( a => n640, b => n641, outb => n639);
   U726 : nand2 port map( a => n643, b => n644, outb => n642);
   U727 : nor2 port map( a => mult_125_G4_ab_4_5_port, b => n646, outb => n645)
                           ;
   U728 : nor2 port map( a => mult_125_G4_ab_5_5_port, b => n648, outb => n647)
                           ;
   U729 : nand2 port map( a => n650, b => n651, outb => n649);
   U730 : nor2 port map( a => mult_125_G4_ab_7_5_port, b => n653, outb => n652)
                           ;
   U731 : nor2 port map( a => mult_125_G4_ab_8_5_port, b => n655, outb => n654)
                           ;
   U732 : nor2 port map( a => mult_125_G4_ab_9_5_port, b => n657, outb => n656)
                           ;
   U733 : nor2 port map( a => mult_125_G4_ab_10_5_port, b => n659, outb => n658
                           );
   U734 : nor2 port map( a => mult_125_G4_ab_11_5_port, b => n661, outb => n660
                           );
   U735 : nor2 port map( a => mult_125_G4_ab_12_5_port, b => n663, outb => n662
                           );
   U736 : nor2 port map( a => mult_125_G4_ab_13_5_port, b => n665, outb => n664
                           );
   U737 : nor2 port map( a => mult_125_G4_ab_14_5_port, b => n667, outb => n666
                           );
   U738 : nand2 port map( a => n669, b => n670, outb => n668);
   U739 : nand2 port map( a => n672, b => n673, outb => n671);
   U740 : nor2 port map( a => mult_125_G4_ab_3_4_port, b => n675, outb => n674)
                           ;
   U741 : nor2 port map( a => mult_125_G4_ab_4_4_port, b => n677, outb => n676)
                           ;
   U742 : nand2 port map( a => n679, b => n680, outb => n678);
   U743 : nor2 port map( a => mult_125_G4_ab_6_4_port, b => n682, outb => n681)
                           ;
   U744 : nand2 port map( a => n684, b => n685, outb => n683);
   U745 : nor2 port map( a => mult_125_G4_ab_8_4_port, b => n687, outb => n686)
                           ;
   U746 : nor2 port map( a => mult_125_G4_ab_9_4_port, b => n689, outb => n688)
                           ;
   U747 : nor2 port map( a => mult_125_G4_ab_10_4_port, b => n691, outb => n690
                           );
   U748 : nand2 port map( a => n693, b => n694, outb => n692);
   U749 : nor2 port map( a => mult_125_G4_ab_12_4_port, b => n696, outb => n695
                           );
   U750 : nor2 port map( a => mult_125_G4_ab_13_4_port, b => n698, outb => n697
                           );
   U751 : nor2 port map( a => mult_125_G4_ab_14_4_port, b => n700, outb => n699
                           );
   U752 : nand2 port map( a => n702, b => n703, outb => n701);
   U753 : nand2 port map( a => n705, b => n706, outb => n704);
   U754 : nand2 port map( a => n708, b => n709, outb => n707);
   U755 : nor2 port map( a => mult_125_G4_ab_4_3_port, b => n711, outb => n710)
                           ;
   U756 : nor2 port map( a => mult_125_G4_ab_5_3_port, b => n713, outb => n712)
                           ;
   U757 : nor2 port map( a => mult_125_G4_ab_6_3_port, b => n715, outb => n714)
                           ;
   U758 : nor2 port map( a => mult_125_G4_ab_7_3_port, b => n717, outb => n716)
                           ;
   U759 : nor2 port map( a => mult_125_G4_ab_8_3_port, b => n719, outb => n718)
                           ;
   U760 : nor2 port map( a => mult_125_G4_ab_9_3_port, b => n721, outb => n720)
                           ;
   U761 : nor2 port map( a => mult_125_G4_ab_10_3_port, b => n723, outb => n722
                           );
   U762 : nor2 port map( a => mult_125_G4_ab_11_3_port, b => n725, outb => n724
                           );
   U763 : nor2 port map( a => mult_125_G4_ab_12_3_port, b => n727, outb => n726
                           );
   U764 : nor2 port map( a => mult_125_G4_ab_13_3_port, b => n729, outb => n728
                           );
   U765 : nor2 port map( a => mult_125_G4_ab_14_3_port, b => n731, outb => n730
                           );
   U766 : nor2 port map( a => mult_125_G4_ab_15_3_port, b => n733, outb => n732
                           );
   U767 : nand2 port map( a => n735, b => n736, outb => n734);
   U768 : nor2 port map( a => mult_125_G4_ab_3_2_port, b => n738, outb => n737)
                           ;
   U769 : nor2 port map( a => mult_125_G4_ab_4_2_port, b => n740, outb => n739)
                           ;
   U770 : nor2 port map( a => mult_125_G4_ab_5_2_port, b => n742, outb => n741)
                           ;
   U771 : nor2 port map( a => mult_125_G4_ab_6_2_port, b => n744, outb => n743)
                           ;
   U772 : nand2 port map( a => n746, b => n747, outb => n745);
   U773 : nor2 port map( a => mult_125_G4_ab_8_2_port, b => n749, outb => n748)
                           ;
   U774 : nor2 port map( a => mult_125_G4_ab_9_2_port, b => n751, outb => n750)
                           ;
   U775 : nor2 port map( a => mult_125_G4_ab_10_2_port, b => n753, outb => n752
                           );
   U776 : nor2 port map( a => mult_125_G4_ab_11_2_port, b => n755, outb => n754
                           );
   U777 : nor2 port map( a => mult_125_G4_ab_12_2_port, b => n757, outb => n756
                           );
   U778 : nor2 port map( a => mult_125_G4_ab_13_2_port, b => n759, outb => n758
                           );
   U779 : nor2 port map( a => mult_125_G4_ab_14_2_port, b => n761, outb => n760
                           );
   U780 : nor2 port map( a => mult_125_G4_ab_15_2_port, b => n763, outb => n762
                           );
   U781 : nand2 port map( a => n765, b => n766, outb => n764);
   U782 : nor2 port map( a => mult_125_G4_ab_3_1_port, b => n768, outb => n767)
                           ;
   U783 : nor2 port map( a => mult_125_G4_ab_4_1_port, b => n770, outb => n769)
                           ;
   U784 : nor2 port map( a => mult_125_G4_ab_5_1_port, b => n772, outb => n771)
                           ;
   U785 : nor2 port map( a => mult_125_G4_ab_6_1_port, b => n774, outb => n773)
                           ;
   U786 : nor2 port map( a => mult_125_G4_ab_7_1_port, b => n776, outb => n775)
                           ;
   U787 : nor2 port map( a => mult_125_G4_ab_8_1_port, b => n778, outb => n777)
                           ;
   U788 : nor2 port map( a => mult_125_G4_ab_9_1_port, b => n780, outb => n779)
                           ;
   U789 : nor2 port map( a => mult_125_G4_ab_10_1_port, b => n782, outb => n781
                           );
   U790 : nor2 port map( a => mult_125_G4_ab_11_1_port, b => n784, outb => n783
                           );
   U791 : nor2 port map( a => mult_125_G4_ab_12_1_port, b => n786, outb => n785
                           );
   U792 : nor2 port map( a => mult_125_G4_ab_13_1_port, b => n788, outb => n787
                           );
   U793 : nor2 port map( a => mult_125_G4_ab_14_1_port, b => n790, outb => n789
                           );
   U794 : nor2 port map( a => mult_125_G4_ab_15_1_port, b => n792, outb => n791
                           );
   U795 : nor2 port map( a => mult_125_G4_ab_2_0_port, b => n794, outb => n793)
                           ;
   U796 : nor2 port map( a => mult_125_G4_ab_3_0_port, b => n796, outb => n795)
                           ;
   U797 : nor2 port map( a => mult_125_G4_ab_4_0_port, b => n798, outb => n797)
                           ;
   U798 : nor2 port map( a => mult_125_G4_ab_5_0_port, b => n800, outb => n799)
                           ;
   U799 : nor2 port map( a => mult_125_G4_ab_6_0_port, b => n802, outb => n801)
                           ;
   U800 : nor2 port map( a => mult_125_G4_ab_7_0_port, b => n804, outb => n803)
                           ;
   U801 : nor2 port map( a => mult_125_G4_ab_8_0_port, b => n806, outb => n805)
                           ;
   U802 : nor2 port map( a => mult_125_G4_ab_9_0_port, b => n808, outb => n807)
                           ;
   U803 : nor2 port map( a => mult_125_G4_ab_10_0_port, b => n810, outb => n809
                           );
   U804 : nor2 port map( a => mult_125_G4_ab_11_0_port, b => n812, outb => n811
                           );
   U805 : nor2 port map( a => mult_125_G4_ab_12_0_port, b => n814, outb => n813
                           );
   U806 : nor2 port map( a => mult_125_G4_ab_13_0_port, b => n816, outb => n815
                           );
   U807 : nor2 port map( a => mult_125_G4_ab_14_0_port, b => n818, outb => n817
                           );
   U808 : nor2 port map( a => mult_125_G4_ab_15_0_port, b => n820, outb => n819
                           );
   U809 : nor2 port map( a => mult_125_G4_ZB, b => mult_125_G4_ZA, outb => n274
                           );
   U810 : nand2 port map( a => mult_125_G4_QB, b => mult_125_G4_ab_15_15_port, 
                           outb => n821);
   U811 : nor2 port map( a => mult_125_G3_ab_1_15_port, b => 
                           mult_125_G3_ab_2_14_port, outb => n822);
   U812 : nor2 port map( a => mult_125_G3_ab_2_15_port, b => 
                           mult_125_G3_ab_3_14_port, outb => n823);
   U813 : nor2 port map( a => mult_125_G3_ab_3_15_port, b => 
                           mult_125_G3_ab_4_14_port, outb => n824);
   U814 : nor2 port map( a => mult_125_G3_ab_4_15_port, b => 
                           mult_125_G3_ab_5_14_port, outb => n825);
   U815 : nor2 port map( a => mult_125_G3_ab_5_15_port, b => 
                           mult_125_G3_ab_6_14_port, outb => n826);
   U816 : nor2 port map( a => mult_125_G3_ab_6_15_port, b => 
                           mult_125_G3_ab_7_14_port, outb => n827);
   U817 : nor2 port map( a => mult_125_G3_ab_7_15_port, b => 
                           mult_125_G3_ab_8_14_port, outb => n828);
   U818 : nor2 port map( a => mult_125_G3_ab_8_15_port, b => 
                           mult_125_G3_ab_9_14_port, outb => n829);
   U819 : nor2 port map( a => mult_125_G3_ab_9_15_port, b => 
                           mult_125_G3_ab_10_14_port, outb => n830);
   U820 : nor2 port map( a => mult_125_G3_ab_10_15_port, b => 
                           mult_125_G3_ab_11_14_port, outb => n831);
   U821 : nor2 port map( a => mult_125_G3_ab_11_15_port, b => 
                           mult_125_G3_ab_12_14_port, outb => n832);
   U822 : nor2 port map( a => mult_125_G3_ab_12_15_port, b => 
                           mult_125_G3_ab_13_14_port, outb => n833);
   U823 : nor2 port map( a => mult_125_G3_ab_13_15_port, b => 
                           mult_125_G3_ab_14_14_port, outb => n834);
   U824 : nor2 port map( a => mult_125_G3_ab_14_15_port, b => 
                           mult_125_G3_ab_15_14_port, outb => n835);
   U825 : nand2 port map( a => n837, b => n838, outb => n836);
   U826 : nand2 port map( a => n840, b => n841, outb => n839);
   U827 : nor2 port map( a => mult_125_G3_ab_4_13_port, b => n843, outb => n842
                           );
   U828 : nor2 port map( a => mult_125_G3_ab_5_13_port, b => n845, outb => n844
                           );
   U829 : nor2 port map( a => mult_125_G3_ab_6_13_port, b => n847, outb => n846
                           );
   U830 : nor2 port map( a => mult_125_G3_ab_7_13_port, b => n849, outb => n848
                           );
   U831 : nor2 port map( a => mult_125_G3_ab_8_13_port, b => n851, outb => n850
                           );
   U832 : nor2 port map( a => mult_125_G3_ab_9_13_port, b => n853, outb => n852
                           );
   U833 : nor2 port map( a => mult_125_G3_ab_10_13_port, b => n855, outb => 
                           n854);
   U834 : nor2 port map( a => mult_125_G3_ab_11_13_port, b => n857, outb => 
                           n856);
   U835 : nor2 port map( a => mult_125_G3_ab_12_13_port, b => n859, outb => 
                           n858);
   U836 : nor2 port map( a => mult_125_G3_ab_13_13_port, b => n861, outb => 
                           n860);
   U837 : nor2 port map( a => mult_125_G3_ab_14_13_port, b => n863, outb => 
                           n862);
   U838 : nor2 port map( a => mult_125_G3_ab_15_13_port, b => n865, outb => 
                           n864);
   U839 : nand2 port map( a => n867, b => n868, outb => n866);
   U840 : nor2 port map( a => mult_125_G3_ab_3_12_port, b => n870, outb => n869
                           );
   U841 : nor2 port map( a => mult_125_G3_ab_4_12_port, b => n872, outb => n871
                           );
   U842 : nor2 port map( a => mult_125_G3_ab_5_12_port, b => n874, outb => n873
                           );
   U843 : nor2 port map( a => mult_125_G3_ab_6_12_port, b => n876, outb => n875
                           );
   U844 : nor2 port map( a => mult_125_G3_ab_7_12_port, b => n878, outb => n877
                           );
   U845 : nor2 port map( a => mult_125_G3_ab_8_12_port, b => n880, outb => n879
                           );
   U846 : nor2 port map( a => mult_125_G3_ab_9_12_port, b => n882, outb => n881
                           );
   U847 : nor2 port map( a => mult_125_G3_ab_10_12_port, b => n884, outb => 
                           n883);
   U848 : nor2 port map( a => mult_125_G3_ab_11_12_port, b => n886, outb => 
                           n885);
   U849 : nor2 port map( a => mult_125_G3_ab_12_12_port, b => n888, outb => 
                           n887);
   U850 : nor2 port map( a => mult_125_G3_ab_13_12_port, b => n890, outb => 
                           n889);
   U851 : nor2 port map( a => mult_125_G3_ab_14_12_port, b => n892, outb => 
                           n891);
   U852 : nor2 port map( a => mult_125_G3_ab_15_12_port, b => n894, outb => 
                           n893);
   U853 : nand2 port map( a => n896, b => n897, outb => n895);
   U854 : nand2 port map( a => n899, b => n900, outb => n898);
   U855 : nor2 port map( a => mult_125_G3_ab_4_11_port, b => n902, outb => n901
                           );
   U856 : nor2 port map( a => mult_125_G3_ab_5_11_port, b => n904, outb => n903
                           );
   U857 : nor2 port map( a => mult_125_G3_ab_6_11_port, b => n906, outb => n905
                           );
   U858 : nor2 port map( a => mult_125_G3_ab_7_11_port, b => n908, outb => n907
                           );
   U859 : nor2 port map( a => mult_125_G3_ab_8_11_port, b => n910, outb => n909
                           );
   U860 : nor2 port map( a => mult_125_G3_ab_9_11_port, b => n912, outb => n911
                           );
   U861 : nor2 port map( a => mult_125_G3_ab_10_11_port, b => n914, outb => 
                           n913);
   U862 : nor2 port map( a => mult_125_G3_ab_11_11_port, b => n916, outb => 
                           n915);
   U863 : nor2 port map( a => mult_125_G3_ab_12_11_port, b => n918, outb => 
                           n917);
   U864 : nor2 port map( a => mult_125_G3_ab_13_11_port, b => n920, outb => 
                           n919);
   U865 : nor2 port map( a => mult_125_G3_ab_14_11_port, b => n922, outb => 
                           n921);
   U866 : nand2 port map( a => n924, b => n925, outb => n923);
   U867 : nand2 port map( a => n927, b => n928, outb => n926);
   U868 : nor2 port map( a => mult_125_G3_ab_3_10_port, b => n930, outb => n929
                           );
   U869 : nor2 port map( a => mult_125_G3_ab_4_10_port, b => n932, outb => n931
                           );
   U870 : nand2 port map( a => n934, b => n935, outb => n933);
   U871 : nor2 port map( a => mult_125_G3_ab_6_10_port, b => n937, outb => n936
                           );
   U872 : nor2 port map( a => mult_125_G3_ab_7_10_port, b => n939, outb => n938
                           );
   U873 : nor2 port map( a => mult_125_G3_ab_8_10_port, b => n941, outb => n940
                           );
   U874 : nor2 port map( a => mult_125_G3_ab_9_10_port, b => n943, outb => n942
                           );
   U875 : nor2 port map( a => mult_125_G3_ab_10_10_port, b => n945, outb => 
                           n944);
   U876 : nor2 port map( a => mult_125_G3_ab_11_10_port, b => n947, outb => 
                           n946);
   U877 : nor2 port map( a => mult_125_G3_ab_12_10_port, b => n949, outb => 
                           n948);
   U878 : nor2 port map( a => mult_125_G3_ab_13_10_port, b => n951, outb => 
                           n950);
   U879 : nor2 port map( a => mult_125_G3_ab_14_10_port, b => n953, outb => 
                           n952);
   U880 : nor2 port map( a => mult_125_G3_ab_15_10_port, b => n955, outb => 
                           n954);
   U881 : nand2 port map( a => n957, b => n958, outb => n956);
   U882 : nor2 port map( a => mult_125_G3_ab_3_9_port, b => n960, outb => n959)
                           ;
   U883 : nor2 port map( a => mult_125_G3_ab_4_9_port, b => n962, outb => n961)
                           ;
   U884 : nor2 port map( a => mult_125_G3_ab_5_9_port, b => n964, outb => n963)
                           ;
   U885 : nor2 port map( a => mult_125_G3_ab_6_9_port, b => n966, outb => n965)
                           ;
   U886 : nor2 port map( a => mult_125_G3_ab_7_9_port, b => n968, outb => n967)
                           ;
   U887 : nor2 port map( a => mult_125_G3_ab_8_9_port, b => n970, outb => n969)
                           ;
   U888 : nor2 port map( a => mult_125_G3_ab_9_9_port, b => n972, outb => n971)
                           ;
   U889 : nor2 port map( a => mult_125_G3_ab_10_9_port, b => n974, outb => n973
                           );
   U890 : nor2 port map( a => mult_125_G3_ab_11_9_port, b => n976, outb => n975
                           );
   U891 : nor2 port map( a => mult_125_G3_ab_12_9_port, b => n978, outb => n977
                           );
   U892 : nor2 port map( a => mult_125_G3_ab_13_9_port, b => n980, outb => n979
                           );
   U893 : nor2 port map( a => mult_125_G3_ab_14_9_port, b => n982, outb => n981
                           );
   U894 : nand2 port map( a => n984, b => n985, outb => n983);
   U895 : nand2 port map( a => n987, b => n988, outb => n986);
   U896 : nor2 port map( a => mult_125_G3_ab_3_8_port, b => n990, outb => n989)
                           ;
   U897 : nor2 port map( a => mult_125_G3_ab_4_8_port, b => n992, outb => n991)
                           ;
   U898 : nor2 port map( a => mult_125_G3_ab_5_8_port, b => n994, outb => n993)
                           ;
   U899 : nor2 port map( a => mult_125_G3_ab_6_8_port, b => n996, outb => n995)
                           ;
   U900 : nor2 port map( a => mult_125_G3_ab_7_8_port, b => n998, outb => n997)
                           ;
   U901 : nor2 port map( a => mult_125_G3_ab_8_8_port, b => n1000, outb => n999
                           );
   U902 : nor2 port map( a => mult_125_G3_ab_9_8_port, b => n1002, outb => 
                           n1001);
   U903 : nor2 port map( a => mult_125_G3_ab_10_8_port, b => n1004, outb => 
                           n1003);
   U904 : nor2 port map( a => mult_125_G3_ab_11_8_port, b => n1006, outb => 
                           n1005);
   U905 : nor2 port map( a => mult_125_G3_ab_12_8_port, b => n1008, outb => 
                           n1007);
   U906 : nor2 port map( a => mult_125_G3_ab_13_8_port, b => n1010, outb => 
                           n1009);
   U907 : nor2 port map( a => mult_125_G3_ab_14_8_port, b => n1012, outb => 
                           n1011);
   U908 : nor2 port map( a => mult_125_G3_ab_15_8_port, b => n1014, outb => 
                           n1013);
   U909 : nand2 port map( a => n1016, b => n1017, outb => n1015);
   U910 : nand2 port map( a => n1019, b => n1020, outb => n1018);
   U911 : nor2 port map( a => mult_125_G3_ab_4_7_port, b => n1022, outb => 
                           n1021);
   U912 : nor2 port map( a => mult_125_G3_ab_5_7_port, b => n1024, outb => 
                           n1023);
   U913 : nor2 port map( a => mult_125_G3_ab_6_7_port, b => n1026, outb => 
                           n1025);
   U914 : nor2 port map( a => mult_125_G3_ab_7_7_port, b => n1028, outb => 
                           n1027);
   U915 : nor2 port map( a => mult_125_G3_ab_8_7_port, b => n1030, outb => 
                           n1029);
   U916 : nor2 port map( a => mult_125_G3_ab_9_7_port, b => n1032, outb => 
                           n1031);
   U917 : nor2 port map( a => mult_125_G3_ab_10_7_port, b => n1034, outb => 
                           n1033);
   U918 : nor2 port map( a => mult_125_G3_ab_11_7_port, b => n1036, outb => 
                           n1035);
   U919 : nor2 port map( a => mult_125_G3_ab_12_7_port, b => n1038, outb => 
                           n1037);
   U920 : nor2 port map( a => mult_125_G3_ab_13_7_port, b => n1040, outb => 
                           n1039);
   U921 : nor2 port map( a => mult_125_G3_ab_14_7_port, b => n1042, outb => 
                           n1041);
   U922 : nand2 port map( a => n1044, b => n1045, outb => n1043);
   U923 : nand2 port map( a => n1047, b => n1048, outb => n1046);
   U924 : nor2 port map( a => mult_125_G3_ab_3_6_port, b => n1050, outb => 
                           n1049);
   U925 : nor2 port map( a => mult_125_G3_ab_4_6_port, b => n1052, outb => 
                           n1051);
   U926 : nand2 port map( a => n1054, b => n1055, outb => n1053);
   U927 : nor2 port map( a => mult_125_G3_ab_6_6_port, b => n1057, outb => 
                           n1056);
   U928 : nor2 port map( a => mult_125_G3_ab_7_6_port, b => n1059, outb => 
                           n1058);
   U929 : nor2 port map( a => mult_125_G3_ab_8_6_port, b => n1061, outb => 
                           n1060);
   U930 : nand2 port map( a => n1063, b => n1064, outb => n1062);
   U931 : nor2 port map( a => mult_125_G3_ab_10_6_port, b => n1066, outb => 
                           n1065);
   U932 : nor2 port map( a => mult_125_G3_ab_11_6_port, b => n1068, outb => 
                           n1067);
   U933 : nor2 port map( a => mult_125_G3_ab_12_6_port, b => n1070, outb => 
                           n1069);
   U934 : nor2 port map( a => mult_125_G3_ab_13_6_port, b => n1072, outb => 
                           n1071);
   U935 : nor2 port map( a => mult_125_G3_ab_14_6_port, b => n1074, outb => 
                           n1073);
   U936 : nor2 port map( a => mult_125_G3_ab_15_6_port, b => n1076, outb => 
                           n1075);
   U937 : nand2 port map( a => n1078, b => n1079, outb => n1077);
   U938 : nand2 port map( a => n1081, b => n1082, outb => n1080);
   U939 : nor2 port map( a => mult_125_G3_ab_4_5_port, b => n1084, outb => 
                           n1083);
   U940 : nor2 port map( a => mult_125_G3_ab_5_5_port, b => n1086, outb => 
                           n1085);
   U941 : nand2 port map( a => n1088, b => n1089, outb => n1087);
   U942 : nor2 port map( a => mult_125_G3_ab_7_5_port, b => n1091, outb => 
                           n1090);
   U943 : nor2 port map( a => mult_125_G3_ab_8_5_port, b => n1093, outb => 
                           n1092);
   U944 : nor2 port map( a => mult_125_G3_ab_9_5_port, b => n1095, outb => 
                           n1094);
   U945 : nor2 port map( a => mult_125_G3_ab_10_5_port, b => n1097, outb => 
                           n1096);
   U946 : nor2 port map( a => mult_125_G3_ab_11_5_port, b => n1099, outb => 
                           n1098);
   U947 : nor2 port map( a => mult_125_G3_ab_12_5_port, b => n1101, outb => 
                           n1100);
   U948 : nor2 port map( a => mult_125_G3_ab_13_5_port, b => n1103, outb => 
                           n1102);
   U949 : nor2 port map( a => mult_125_G3_ab_14_5_port, b => n1105, outb => 
                           n1104);
   U950 : nand2 port map( a => n1107, b => n1108, outb => n1106);
   U951 : nand2 port map( a => n1110, b => n1111, outb => n1109);
   U952 : nor2 port map( a => mult_125_G3_ab_3_4_port, b => n1113, outb => 
                           n1112);
   U953 : nor2 port map( a => mult_125_G3_ab_4_4_port, b => n1115, outb => 
                           n1114);
   U954 : nand2 port map( a => n1117, b => n1118, outb => n1116);
   U955 : nor2 port map( a => mult_125_G3_ab_6_4_port, b => n1120, outb => 
                           n1119);
   U956 : nand2 port map( a => n1122, b => n1123, outb => n1121);
   U957 : nor2 port map( a => mult_125_G3_ab_8_4_port, b => n1125, outb => 
                           n1124);
   U958 : nor2 port map( a => mult_125_G3_ab_9_4_port, b => n1127, outb => 
                           n1126);
   U959 : nor2 port map( a => mult_125_G3_ab_10_4_port, b => n1129, outb => 
                           n1128);
   U960 : nand2 port map( a => n1131, b => n1132, outb => n1130);
   U961 : nor2 port map( a => mult_125_G3_ab_12_4_port, b => n1134, outb => 
                           n1133);
   U962 : nor2 port map( a => mult_125_G3_ab_13_4_port, b => n1136, outb => 
                           n1135);
   U963 : nor2 port map( a => mult_125_G3_ab_14_4_port, b => n1138, outb => 
                           n1137);
   U964 : nand2 port map( a => n1140, b => n1141, outb => n1139);
   U965 : nand2 port map( a => n1143, b => n1144, outb => n1142);
   U966 : nand2 port map( a => n1146, b => n1147, outb => n1145);
   U967 : nor2 port map( a => mult_125_G3_ab_4_3_port, b => n1149, outb => 
                           n1148);
   U968 : nor2 port map( a => mult_125_G3_ab_5_3_port, b => n1151, outb => 
                           n1150);
   U969 : nor2 port map( a => mult_125_G3_ab_6_3_port, b => n1153, outb => 
                           n1152);
   U970 : nor2 port map( a => mult_125_G3_ab_7_3_port, b => n1155, outb => 
                           n1154);
   U971 : nor2 port map( a => mult_125_G3_ab_8_3_port, b => n1157, outb => 
                           n1156);
   U972 : nor2 port map( a => mult_125_G3_ab_9_3_port, b => n1159, outb => 
                           n1158);
   U973 : nor2 port map( a => mult_125_G3_ab_10_3_port, b => n1161, outb => 
                           n1160);
   U974 : nor2 port map( a => mult_125_G3_ab_11_3_port, b => n1163, outb => 
                           n1162);
   U975 : nor2 port map( a => mult_125_G3_ab_12_3_port, b => n1165, outb => 
                           n1164);
   U976 : nor2 port map( a => mult_125_G3_ab_13_3_port, b => n1167, outb => 
                           n1166);
   U977 : nor2 port map( a => mult_125_G3_ab_14_3_port, b => n1169, outb => 
                           n1168);
   U978 : nor2 port map( a => mult_125_G3_ab_15_3_port, b => n1171, outb => 
                           n1170);
   U979 : nand2 port map( a => n1173, b => n1174, outb => n1172);
   U980 : nor2 port map( a => mult_125_G3_ab_3_2_port, b => n1176, outb => 
                           n1175);
   U981 : nor2 port map( a => mult_125_G3_ab_4_2_port, b => n1178, outb => 
                           n1177);
   U982 : nor2 port map( a => mult_125_G3_ab_5_2_port, b => n1180, outb => 
                           n1179);
   U983 : nor2 port map( a => mult_125_G3_ab_6_2_port, b => n1182, outb => 
                           n1181);
   U984 : nand2 port map( a => n1184, b => n1185, outb => n1183);
   U985 : nor2 port map( a => mult_125_G3_ab_8_2_port, b => n1187, outb => 
                           n1186);
   U986 : nor2 port map( a => mult_125_G3_ab_9_2_port, b => n1189, outb => 
                           n1188);
   U987 : nor2 port map( a => mult_125_G3_ab_10_2_port, b => n1191, outb => 
                           n1190);
   U988 : nor2 port map( a => mult_125_G3_ab_11_2_port, b => n1193, outb => 
                           n1192);
   U989 : nor2 port map( a => mult_125_G3_ab_12_2_port, b => n1195, outb => 
                           n1194);
   U990 : nor2 port map( a => mult_125_G3_ab_13_2_port, b => n1197, outb => 
                           n1196);
   U991 : nor2 port map( a => mult_125_G3_ab_14_2_port, b => n1199, outb => 
                           n1198);
   U992 : nor2 port map( a => mult_125_G3_ab_15_2_port, b => n1201, outb => 
                           n1200);
   U993 : nand2 port map( a => n1203, b => n1204, outb => n1202);
   U994 : nor2 port map( a => mult_125_G3_ab_3_1_port, b => n1206, outb => 
                           n1205);
   U995 : nor2 port map( a => mult_125_G3_ab_4_1_port, b => n1208, outb => 
                           n1207);
   U996 : nor2 port map( a => mult_125_G3_ab_5_1_port, b => n1210, outb => 
                           n1209);
   U997 : nor2 port map( a => mult_125_G3_ab_6_1_port, b => n1212, outb => 
                           n1211);
   U998 : nor2 port map( a => mult_125_G3_ab_7_1_port, b => n1214, outb => 
                           n1213);
   U999 : nor2 port map( a => mult_125_G3_ab_8_1_port, b => n1216, outb => 
                           n1215);
   U1000 : nor2 port map( a => mult_125_G3_ab_9_1_port, b => n1218, outb => 
                           n1217);
   U1001 : nor2 port map( a => mult_125_G3_ab_10_1_port, b => n1220, outb => 
                           n1219);
   U1002 : nor2 port map( a => mult_125_G3_ab_11_1_port, b => n1222, outb => 
                           n1221);
   U1003 : nor2 port map( a => mult_125_G3_ab_12_1_port, b => n1224, outb => 
                           n1223);
   U1004 : nor2 port map( a => mult_125_G3_ab_13_1_port, b => n1226, outb => 
                           n1225);
   U1005 : nor2 port map( a => mult_125_G3_ab_14_1_port, b => n1228, outb => 
                           n1227);
   U1006 : nor2 port map( a => mult_125_G3_ab_15_1_port, b => n1230, outb => 
                           n1229);
   U1007 : nor2 port map( a => mult_125_G3_ab_2_0_port, b => n1232, outb => 
                           n1231);
   U1008 : nor2 port map( a => mult_125_G3_ab_3_0_port, b => n1234, outb => 
                           n1233);
   U1009 : nor2 port map( a => mult_125_G3_ab_4_0_port, b => n1236, outb => 
                           n1235);
   U1010 : nor2 port map( a => mult_125_G3_ab_5_0_port, b => n1238, outb => 
                           n1237);
   U1011 : nor2 port map( a => mult_125_G3_ab_6_0_port, b => n1240, outb => 
                           n1239);
   U1012 : nor2 port map( a => mult_125_G3_ab_7_0_port, b => n1242, outb => 
                           n1241);
   U1013 : nor2 port map( a => mult_125_G3_ab_8_0_port, b => n1244, outb => 
                           n1243);
   U1014 : nor2 port map( a => mult_125_G3_ab_9_0_port, b => n1246, outb => 
                           n1245);
   U1015 : nor2 port map( a => mult_125_G3_ab_10_0_port, b => n1248, outb => 
                           n1247);
   U1016 : nor2 port map( a => mult_125_G3_ab_11_0_port, b => n1250, outb => 
                           n1249);
   U1017 : nor2 port map( a => mult_125_G3_ab_12_0_port, b => n1252, outb => 
                           n1251);
   U1018 : nor2 port map( a => mult_125_G3_ab_13_0_port, b => n1254, outb => 
                           n1253);
   U1019 : nor2 port map( a => mult_125_G3_ab_14_0_port, b => n1256, outb => 
                           n1255);
   U1020 : nor2 port map( a => mult_125_G3_ab_15_0_port, b => n1258, outb => 
                           n1257);
   U1021 : nor2 port map( a => mult_125_G3_ZB, b => mult_125_G3_ZA, outb => 
                           n382);
   U1022 : nand2 port map( a => mult_125_G3_QB, b => mult_125_G3_ab_15_15_port,
                           outb => n1259);
   U1023 : nor2 port map( a => mult_125_G2_ab_1_15_port, b => 
                           mult_125_G2_ab_2_14_port, outb => n1260);
   U1024 : nor2 port map( a => mult_125_G2_ab_2_15_port, b => 
                           mult_125_G2_ab_3_14_port, outb => n1261);
   U1025 : nor2 port map( a => mult_125_G2_ab_3_15_port, b => 
                           mult_125_G2_ab_4_14_port, outb => n1262);
   U1026 : nor2 port map( a => mult_125_G2_ab_4_15_port, b => 
                           mult_125_G2_ab_5_14_port, outb => n1263);
   U1027 : nor2 port map( a => mult_125_G2_ab_5_15_port, b => 
                           mult_125_G2_ab_6_14_port, outb => n1264);
   U1028 : nor2 port map( a => mult_125_G2_ab_6_15_port, b => 
                           mult_125_G2_ab_7_14_port, outb => n1265);
   U1029 : nor2 port map( a => mult_125_G2_ab_7_15_port, b => 
                           mult_125_G2_ab_8_14_port, outb => n1266);
   U1030 : nor2 port map( a => mult_125_G2_ab_8_15_port, b => 
                           mult_125_G2_ab_9_14_port, outb => n1267);
   U1031 : nor2 port map( a => mult_125_G2_ab_9_15_port, b => 
                           mult_125_G2_ab_10_14_port, outb => n1268);
   U1032 : nor2 port map( a => mult_125_G2_ab_10_15_port, b => 
                           mult_125_G2_ab_11_14_port, outb => n1269);
   U1033 : nor2 port map( a => mult_125_G2_ab_11_15_port, b => 
                           mult_125_G2_ab_12_14_port, outb => n1270);
   U1034 : nor2 port map( a => mult_125_G2_ab_12_15_port, b => 
                           mult_125_G2_ab_13_14_port, outb => n1271);
   U1035 : nor2 port map( a => mult_125_G2_ab_13_15_port, b => 
                           mult_125_G2_ab_14_14_port, outb => n1272);
   U1036 : nor2 port map( a => mult_125_G2_ab_14_15_port, b => 
                           mult_125_G2_ab_15_14_port, outb => n1273);
   U1037 : nand2 port map( a => n1275, b => n1276, outb => n1274);
   U1038 : nand2 port map( a => n1278, b => n1279, outb => n1277);
   U1039 : nor2 port map( a => mult_125_G2_ab_4_13_port, b => n1281, outb => 
                           n1280);
   U1040 : nor2 port map( a => mult_125_G2_ab_5_13_port, b => n1283, outb => 
                           n1282);
   U1041 : nor2 port map( a => mult_125_G2_ab_6_13_port, b => n1285, outb => 
                           n1284);
   U1042 : nor2 port map( a => mult_125_G2_ab_7_13_port, b => n1287, outb => 
                           n1286);
   U1043 : nor2 port map( a => mult_125_G2_ab_8_13_port, b => n1289, outb => 
                           n1288);
   U1044 : nor2 port map( a => mult_125_G2_ab_9_13_port, b => n1291, outb => 
                           n1290);
   U1045 : nor2 port map( a => mult_125_G2_ab_10_13_port, b => n1293, outb => 
                           n1292);
   U1046 : nor2 port map( a => mult_125_G2_ab_11_13_port, b => n1295, outb => 
                           n1294);
   U1047 : nor2 port map( a => mult_125_G2_ab_12_13_port, b => n1297, outb => 
                           n1296);
   U1048 : nor2 port map( a => mult_125_G2_ab_13_13_port, b => n1299, outb => 
                           n1298);
   U1049 : nor2 port map( a => mult_125_G2_ab_14_13_port, b => n1301, outb => 
                           n1300);
   U1050 : nor2 port map( a => mult_125_G2_ab_15_13_port, b => n1303, outb => 
                           n1302);
   U1051 : nand2 port map( a => n1305, b => n1306, outb => n1304);
   U1052 : nor2 port map( a => mult_125_G2_ab_3_12_port, b => n1308, outb => 
                           n1307);
   U1053 : nor2 port map( a => mult_125_G2_ab_4_12_port, b => n1310, outb => 
                           n1309);
   U1054 : nor2 port map( a => mult_125_G2_ab_5_12_port, b => n1312, outb => 
                           n1311);
   U1055 : nor2 port map( a => mult_125_G2_ab_6_12_port, b => n1314, outb => 
                           n1313);
   U1056 : nor2 port map( a => mult_125_G2_ab_7_12_port, b => n1316, outb => 
                           n1315);
   U1057 : nor2 port map( a => mult_125_G2_ab_8_12_port, b => n1318, outb => 
                           n1317);
   U1058 : nor2 port map( a => mult_125_G2_ab_9_12_port, b => n1320, outb => 
                           n1319);
   U1059 : nor2 port map( a => mult_125_G2_ab_10_12_port, b => n1322, outb => 
                           n1321);
   U1060 : nor2 port map( a => mult_125_G2_ab_11_12_port, b => n1324, outb => 
                           n1323);
   U1061 : nor2 port map( a => mult_125_G2_ab_12_12_port, b => n1326, outb => 
                           n1325);
   U1062 : nor2 port map( a => mult_125_G2_ab_13_12_port, b => n1328, outb => 
                           n1327);
   U1063 : nor2 port map( a => mult_125_G2_ab_14_12_port, b => n1330, outb => 
                           n1329);
   U1064 : nor2 port map( a => mult_125_G2_ab_15_12_port, b => n1332, outb => 
                           n1331);
   U1065 : nand2 port map( a => n1334, b => n1335, outb => n1333);
   U1066 : nand2 port map( a => n1337, b => n1338, outb => n1336);
   U1067 : nor2 port map( a => mult_125_G2_ab_4_11_port, b => n1340, outb => 
                           n1339);
   U1068 : nor2 port map( a => mult_125_G2_ab_5_11_port, b => n1342, outb => 
                           n1341);
   U1069 : nor2 port map( a => mult_125_G2_ab_6_11_port, b => n1344, outb => 
                           n1343);
   U1070 : nor2 port map( a => mult_125_G2_ab_7_11_port, b => n1346, outb => 
                           n1345);
   U1071 : nor2 port map( a => mult_125_G2_ab_8_11_port, b => n1348, outb => 
                           n1347);
   U1072 : nor2 port map( a => mult_125_G2_ab_9_11_port, b => n1350, outb => 
                           n1349);
   U1073 : nor2 port map( a => mult_125_G2_ab_10_11_port, b => n1352, outb => 
                           n1351);
   U1074 : nor2 port map( a => mult_125_G2_ab_11_11_port, b => n1354, outb => 
                           n1353);
   U1075 : nor2 port map( a => mult_125_G2_ab_12_11_port, b => n1356, outb => 
                           n1355);
   U1076 : nor2 port map( a => mult_125_G2_ab_13_11_port, b => n1358, outb => 
                           n1357);
   U1077 : nor2 port map( a => mult_125_G2_ab_14_11_port, b => n1360, outb => 
                           n1359);
   U1078 : nand2 port map( a => n1362, b => n1363, outb => n1361);
   U1079 : nand2 port map( a => n1365, b => n1366, outb => n1364);
   U1080 : nor2 port map( a => mult_125_G2_ab_3_10_port, b => n1368, outb => 
                           n1367);
   U1081 : nor2 port map( a => mult_125_G2_ab_4_10_port, b => n1370, outb => 
                           n1369);
   U1082 : nand2 port map( a => n1372, b => n1373, outb => n1371);
   U1083 : nor2 port map( a => mult_125_G2_ab_6_10_port, b => n1375, outb => 
                           n1374);
   U1084 : nor2 port map( a => mult_125_G2_ab_7_10_port, b => n1377, outb => 
                           n1376);
   U1085 : nor2 port map( a => mult_125_G2_ab_8_10_port, b => n1379, outb => 
                           n1378);
   U1086 : nor2 port map( a => mult_125_G2_ab_9_10_port, b => n1381, outb => 
                           n1380);
   U1087 : nor2 port map( a => mult_125_G2_ab_10_10_port, b => n1383, outb => 
                           n1382);
   U1088 : nor2 port map( a => mult_125_G2_ab_11_10_port, b => n1385, outb => 
                           n1384);
   U1089 : nor2 port map( a => mult_125_G2_ab_12_10_port, b => n1387, outb => 
                           n1386);
   U1090 : nor2 port map( a => mult_125_G2_ab_13_10_port, b => n1389, outb => 
                           n1388);
   U1091 : nor2 port map( a => mult_125_G2_ab_14_10_port, b => n1391, outb => 
                           n1390);
   U1092 : nor2 port map( a => mult_125_G2_ab_15_10_port, b => n1393, outb => 
                           n1392);
   U1093 : nand2 port map( a => n1395, b => n1396, outb => n1394);
   U1094 : nor2 port map( a => mult_125_G2_ab_3_9_port, b => n1398, outb => 
                           n1397);
   U1095 : nor2 port map( a => mult_125_G2_ab_4_9_port, b => n1400, outb => 
                           n1399);
   U1096 : nor2 port map( a => mult_125_G2_ab_5_9_port, b => n1402, outb => 
                           n1401);
   U1097 : nor2 port map( a => mult_125_G2_ab_6_9_port, b => n1404, outb => 
                           n1403);
   U1098 : nor2 port map( a => mult_125_G2_ab_7_9_port, b => n1406, outb => 
                           n1405);
   U1099 : nor2 port map( a => mult_125_G2_ab_8_9_port, b => n1408, outb => 
                           n1407);
   U1100 : nor2 port map( a => mult_125_G2_ab_9_9_port, b => n1410, outb => 
                           n1409);
   U1101 : nor2 port map( a => mult_125_G2_ab_10_9_port, b => n1412, outb => 
                           n1411);
   U1102 : nor2 port map( a => mult_125_G2_ab_11_9_port, b => n1414, outb => 
                           n1413);
   U1103 : nor2 port map( a => mult_125_G2_ab_12_9_port, b => n1416, outb => 
                           n1415);
   U1104 : nor2 port map( a => mult_125_G2_ab_13_9_port, b => n1418, outb => 
                           n1417);
   U1105 : nor2 port map( a => mult_125_G2_ab_14_9_port, b => n1420, outb => 
                           n1419);
   U1106 : nand2 port map( a => n1422, b => n1423, outb => n1421);
   U1107 : nand2 port map( a => n1425, b => n1426, outb => n1424);
   U1108 : nor2 port map( a => mult_125_G2_ab_3_8_port, b => n1428, outb => 
                           n1427);
   U1109 : nor2 port map( a => mult_125_G2_ab_4_8_port, b => n1430, outb => 
                           n1429);
   U1110 : nor2 port map( a => mult_125_G2_ab_5_8_port, b => n1432, outb => 
                           n1431);
   U1111 : nor2 port map( a => mult_125_G2_ab_6_8_port, b => n1434, outb => 
                           n1433);
   U1112 : nor2 port map( a => mult_125_G2_ab_7_8_port, b => n1436, outb => 
                           n1435);
   U1113 : nor2 port map( a => mult_125_G2_ab_8_8_port, b => n1438, outb => 
                           n1437);
   U1114 : nor2 port map( a => mult_125_G2_ab_9_8_port, b => n1440, outb => 
                           n1439);
   U1115 : nor2 port map( a => mult_125_G2_ab_10_8_port, b => n1442, outb => 
                           n1441);
   U1116 : nor2 port map( a => mult_125_G2_ab_11_8_port, b => n1444, outb => 
                           n1443);
   U1117 : nor2 port map( a => mult_125_G2_ab_12_8_port, b => n1446, outb => 
                           n1445);
   U1118 : nor2 port map( a => mult_125_G2_ab_13_8_port, b => n1448, outb => 
                           n1447);
   U1119 : nor2 port map( a => mult_125_G2_ab_14_8_port, b => n1450, outb => 
                           n1449);
   U1120 : nor2 port map( a => mult_125_G2_ab_15_8_port, b => n1452, outb => 
                           n1451);
   U1121 : nand2 port map( a => n1454, b => n1455, outb => n1453);
   U1122 : nand2 port map( a => n1457, b => n1458, outb => n1456);
   U1123 : nor2 port map( a => mult_125_G2_ab_4_7_port, b => n1460, outb => 
                           n1459);
   U1124 : nor2 port map( a => mult_125_G2_ab_5_7_port, b => n1462, outb => 
                           n1461);
   U1125 : nor2 port map( a => mult_125_G2_ab_6_7_port, b => n1464, outb => 
                           n1463);
   U1126 : nor2 port map( a => mult_125_G2_ab_7_7_port, b => n1466, outb => 
                           n1465);
   U1127 : nor2 port map( a => mult_125_G2_ab_8_7_port, b => n1468, outb => 
                           n1467);
   U1128 : nor2 port map( a => mult_125_G2_ab_9_7_port, b => n1470, outb => 
                           n1469);
   U1129 : nor2 port map( a => mult_125_G2_ab_10_7_port, b => n1472, outb => 
                           n1471);
   U1130 : nor2 port map( a => mult_125_G2_ab_11_7_port, b => n1474, outb => 
                           n1473);
   U1131 : nor2 port map( a => mult_125_G2_ab_12_7_port, b => n1476, outb => 
                           n1475);
   U1132 : nor2 port map( a => mult_125_G2_ab_13_7_port, b => n1478, outb => 
                           n1477);
   U1133 : nor2 port map( a => mult_125_G2_ab_14_7_port, b => n1480, outb => 
                           n1479);
   U1134 : nand2 port map( a => n1482, b => n1483, outb => n1481);
   U1135 : nand2 port map( a => n1485, b => n1486, outb => n1484);
   U1136 : nor2 port map( a => mult_125_G2_ab_3_6_port, b => n1488, outb => 
                           n1487);
   U1137 : nor2 port map( a => mult_125_G2_ab_4_6_port, b => n1490, outb => 
                           n1489);
   U1138 : nand2 port map( a => n1492, b => n1493, outb => n1491);
   U1139 : nor2 port map( a => mult_125_G2_ab_6_6_port, b => n1495, outb => 
                           n1494);
   U1140 : nor2 port map( a => mult_125_G2_ab_7_6_port, b => n1497, outb => 
                           n1496);
   U1141 : nor2 port map( a => mult_125_G2_ab_8_6_port, b => n1499, outb => 
                           n1498);
   U1142 : nand2 port map( a => n1501, b => n1502, outb => n1500);
   U1143 : nor2 port map( a => mult_125_G2_ab_10_6_port, b => n1504, outb => 
                           n1503);
   U1144 : nor2 port map( a => mult_125_G2_ab_11_6_port, b => n1506, outb => 
                           n1505);
   U1145 : nor2 port map( a => mult_125_G2_ab_12_6_port, b => n1508, outb => 
                           n1507);
   U1146 : nor2 port map( a => mult_125_G2_ab_13_6_port, b => n1510, outb => 
                           n1509);
   U1147 : nor2 port map( a => mult_125_G2_ab_14_6_port, b => n1512, outb => 
                           n1511);
   U1148 : nor2 port map( a => mult_125_G2_ab_15_6_port, b => n1514, outb => 
                           n1513);
   U1149 : nand2 port map( a => n1516, b => n1517, outb => n1515);
   U1150 : nand2 port map( a => n1519, b => n1520, outb => n1518);
   U1151 : nor2 port map( a => mult_125_G2_ab_4_5_port, b => n1522, outb => 
                           n1521);
   U1152 : nor2 port map( a => mult_125_G2_ab_5_5_port, b => n1524, outb => 
                           n1523);
   U1153 : nand2 port map( a => n1526, b => n1527, outb => n1525);
   U1154 : nor2 port map( a => mult_125_G2_ab_7_5_port, b => n1529, outb => 
                           n1528);
   U1155 : nor2 port map( a => mult_125_G2_ab_8_5_port, b => n1531, outb => 
                           n1530);
   U1156 : nor2 port map( a => mult_125_G2_ab_9_5_port, b => n1533, outb => 
                           n1532);
   U1157 : nor2 port map( a => mult_125_G2_ab_10_5_port, b => n1535, outb => 
                           n1534);
   U1158 : nor2 port map( a => mult_125_G2_ab_11_5_port, b => n1537, outb => 
                           n1536);
   U1159 : nor2 port map( a => mult_125_G2_ab_12_5_port, b => n1539, outb => 
                           n1538);
   U1160 : nor2 port map( a => mult_125_G2_ab_13_5_port, b => n1541, outb => 
                           n1540);
   U1161 : nor2 port map( a => mult_125_G2_ab_14_5_port, b => n1543, outb => 
                           n1542);
   U1162 : nand2 port map( a => n1545, b => n1546, outb => n1544);
   U1163 : nand2 port map( a => n1548, b => n1549, outb => n1547);
   U1164 : nor2 port map( a => mult_125_G2_ab_3_4_port, b => n1551, outb => 
                           n1550);
   U1165 : nor2 port map( a => mult_125_G2_ab_4_4_port, b => n1553, outb => 
                           n1552);
   U1166 : nand2 port map( a => n1555, b => n1556, outb => n1554);
   U1167 : nor2 port map( a => mult_125_G2_ab_6_4_port, b => n1558, outb => 
                           n1557);
   U1168 : nand2 port map( a => n1560, b => n1561, outb => n1559);
   U1169 : nor2 port map( a => mult_125_G2_ab_8_4_port, b => n1563, outb => 
                           n1562);
   U1170 : nor2 port map( a => mult_125_G2_ab_9_4_port, b => n1565, outb => 
                           n1564);
   U1171 : nor2 port map( a => mult_125_G2_ab_10_4_port, b => n1567, outb => 
                           n1566);
   U1172 : nand2 port map( a => n1569, b => n1570, outb => n1568);
   U1173 : nor2 port map( a => mult_125_G2_ab_12_4_port, b => n1572, outb => 
                           n1571);
   U1174 : nor2 port map( a => mult_125_G2_ab_13_4_port, b => n1574, outb => 
                           n1573);
   U1175 : nor2 port map( a => mult_125_G2_ab_14_4_port, b => n1576, outb => 
                           n1575);
   U1176 : nand2 port map( a => n1578, b => n1579, outb => n1577);
   U1177 : nand2 port map( a => n1581, b => n1582, outb => n1580);
   U1178 : nand2 port map( a => n1584, b => n1585, outb => n1583);
   U1179 : nor2 port map( a => mult_125_G2_ab_4_3_port, b => n1587, outb => 
                           n1586);
   U1180 : nor2 port map( a => mult_125_G2_ab_5_3_port, b => n1589, outb => 
                           n1588);
   U1181 : nor2 port map( a => mult_125_G2_ab_6_3_port, b => n1591, outb => 
                           n1590);
   U1182 : nor2 port map( a => mult_125_G2_ab_7_3_port, b => n1593, outb => 
                           n1592);
   U1183 : nor2 port map( a => mult_125_G2_ab_8_3_port, b => n1595, outb => 
                           n1594);
   U1184 : nor2 port map( a => mult_125_G2_ab_9_3_port, b => n1597, outb => 
                           n1596);
   U1185 : nor2 port map( a => mult_125_G2_ab_10_3_port, b => n1599, outb => 
                           n1598);
   U1186 : nor2 port map( a => mult_125_G2_ab_11_3_port, b => n1601, outb => 
                           n1600);
   U1187 : nor2 port map( a => mult_125_G2_ab_12_3_port, b => n1603, outb => 
                           n1602);
   U1188 : nor2 port map( a => mult_125_G2_ab_13_3_port, b => n1605, outb => 
                           n1604);
   U1189 : nor2 port map( a => mult_125_G2_ab_14_3_port, b => n1607, outb => 
                           n1606);
   U1190 : nor2 port map( a => mult_125_G2_ab_15_3_port, b => n1609, outb => 
                           n1608);
   U1191 : nand2 port map( a => n1611, b => n1612, outb => n1610);
   U1192 : nor2 port map( a => mult_125_G2_ab_3_2_port, b => n1614, outb => 
                           n1613);
   U1193 : nor2 port map( a => mult_125_G2_ab_4_2_port, b => n1616, outb => 
                           n1615);
   U1194 : nor2 port map( a => mult_125_G2_ab_5_2_port, b => n1618, outb => 
                           n1617);
   U1195 : nor2 port map( a => mult_125_G2_ab_6_2_port, b => n1620, outb => 
                           n1619);
   U1196 : nand2 port map( a => n1622, b => n1623, outb => n1621);
   U1197 : nor2 port map( a => mult_125_G2_ab_8_2_port, b => n1625, outb => 
                           n1624);
   U1198 : nor2 port map( a => mult_125_G2_ab_9_2_port, b => n1627, outb => 
                           n1626);
   U1199 : nor2 port map( a => mult_125_G2_ab_10_2_port, b => n1629, outb => 
                           n1628);
   U1200 : nor2 port map( a => mult_125_G2_ab_11_2_port, b => n1631, outb => 
                           n1630);
   U1201 : nor2 port map( a => mult_125_G2_ab_12_2_port, b => n1633, outb => 
                           n1632);
   U1202 : nor2 port map( a => mult_125_G2_ab_13_2_port, b => n1635, outb => 
                           n1634);
   U1203 : nor2 port map( a => mult_125_G2_ab_14_2_port, b => n1637, outb => 
                           n1636);
   U1204 : nor2 port map( a => mult_125_G2_ab_15_2_port, b => n1639, outb => 
                           n1638);
   U1205 : nand2 port map( a => n1641, b => n1642, outb => n1640);
   U1206 : nor2 port map( a => mult_125_G2_ab_3_1_port, b => n1644, outb => 
                           n1643);
   U1207 : nor2 port map( a => mult_125_G2_ab_4_1_port, b => n1646, outb => 
                           n1645);
   U1208 : nor2 port map( a => mult_125_G2_ab_5_1_port, b => n1648, outb => 
                           n1647);
   U1209 : nor2 port map( a => mult_125_G2_ab_6_1_port, b => n1650, outb => 
                           n1649);
   U1210 : nor2 port map( a => mult_125_G2_ab_7_1_port, b => n1652, outb => 
                           n1651);
   U1211 : nor2 port map( a => mult_125_G2_ab_8_1_port, b => n1654, outb => 
                           n1653);
   U1212 : nor2 port map( a => mult_125_G2_ab_9_1_port, b => n1656, outb => 
                           n1655);
   U1213 : nor2 port map( a => mult_125_G2_ab_10_1_port, b => n1658, outb => 
                           n1657);
   U1214 : nor2 port map( a => mult_125_G2_ab_11_1_port, b => n1660, outb => 
                           n1659);
   U1215 : nor2 port map( a => mult_125_G2_ab_12_1_port, b => n1662, outb => 
                           n1661);
   U1216 : nor2 port map( a => mult_125_G2_ab_13_1_port, b => n1664, outb => 
                           n1663);
   U1217 : nor2 port map( a => mult_125_G2_ab_14_1_port, b => n1666, outb => 
                           n1665);
   U1218 : nor2 port map( a => mult_125_G2_ab_15_1_port, b => n1668, outb => 
                           n1667);
   U1219 : nor2 port map( a => mult_125_G2_ab_2_0_port, b => n1670, outb => 
                           n1669);
   U1220 : nor2 port map( a => mult_125_G2_ab_3_0_port, b => n1672, outb => 
                           n1671);
   U1221 : nor2 port map( a => mult_125_G2_ab_4_0_port, b => n1674, outb => 
                           n1673);
   U1222 : nor2 port map( a => mult_125_G2_ab_5_0_port, b => n1676, outb => 
                           n1675);
   U1223 : nor2 port map( a => mult_125_G2_ab_6_0_port, b => n1678, outb => 
                           n1677);
   U1224 : nor2 port map( a => mult_125_G2_ab_7_0_port, b => n1680, outb => 
                           n1679);
   U1225 : nor2 port map( a => mult_125_G2_ab_8_0_port, b => n1682, outb => 
                           n1681);
   U1226 : nor2 port map( a => mult_125_G2_ab_9_0_port, b => n1684, outb => 
                           n1683);
   U1227 : nor2 port map( a => mult_125_G2_ab_10_0_port, b => n1686, outb => 
                           n1685);
   U1228 : nor2 port map( a => mult_125_G2_ab_11_0_port, b => n1688, outb => 
                           n1687);
   U1229 : nor2 port map( a => mult_125_G2_ab_12_0_port, b => n1690, outb => 
                           n1689);
   U1230 : nor2 port map( a => mult_125_G2_ab_13_0_port, b => n1692, outb => 
                           n1691);
   U1231 : nor2 port map( a => mult_125_G2_ab_14_0_port, b => n1694, outb => 
                           n1693);
   U1232 : nor2 port map( a => mult_125_G2_ab_15_0_port, b => n1696, outb => 
                           n1695);
   U1233 : nor2 port map( a => mult_125_G2_ZB, b => mult_125_G2_ZA, outb => 
                           n346);
   U1234 : nand2 port map( a => mult_125_G2_QB, b => mult_125_G2_ab_15_15_port,
                           outb => n1697);
   U1235 : nor2 port map( a => mult_125_ab_1_15_port, b => 
                           mult_125_ab_2_14_port, outb => n1698);
   U1236 : nor2 port map( a => mult_125_ab_2_15_port, b => 
                           mult_125_ab_3_14_port, outb => n1699);
   U1237 : nor2 port map( a => mult_125_ab_3_15_port, b => 
                           mult_125_ab_4_14_port, outb => n1700);
   U1238 : nor2 port map( a => mult_125_ab_4_15_port, b => 
                           mult_125_ab_5_14_port, outb => n1701);
   U1239 : nor2 port map( a => mult_125_ab_5_15_port, b => 
                           mult_125_ab_6_14_port, outb => n1702);
   U1240 : nor2 port map( a => mult_125_ab_6_15_port, b => 
                           mult_125_ab_7_14_port, outb => n1703);
   U1241 : nor2 port map( a => mult_125_ab_7_15_port, b => 
                           mult_125_ab_8_14_port, outb => n1704);
   U1242 : nor2 port map( a => mult_125_ab_8_15_port, b => 
                           mult_125_ab_9_14_port, outb => n1705);
   U1243 : nor2 port map( a => mult_125_ab_9_15_port, b => 
                           mult_125_ab_10_14_port, outb => n1706);
   U1244 : nor2 port map( a => mult_125_ab_10_15_port, b => 
                           mult_125_ab_11_14_port, outb => n1707);
   U1245 : nor2 port map( a => mult_125_ab_11_15_port, b => 
                           mult_125_ab_12_14_port, outb => n1708);
   U1246 : nor2 port map( a => mult_125_ab_12_15_port, b => 
                           mult_125_ab_13_14_port, outb => n1709);
   U1247 : nor2 port map( a => mult_125_ab_13_15_port, b => 
                           mult_125_ab_14_14_port, outb => n1710);
   U1248 : nor2 port map( a => mult_125_ab_14_15_port, b => 
                           mult_125_ab_15_14_port, outb => n1711);
   U1249 : nand2 port map( a => n1713, b => n1714, outb => n1712);
   U1250 : nand2 port map( a => n1716, b => n1717, outb => n1715);
   U1251 : nor2 port map( a => mult_125_ab_4_13_port, b => n1719, outb => n1718
                           );
   U1252 : nor2 port map( a => mult_125_ab_5_13_port, b => n1721, outb => n1720
                           );
   U1253 : nor2 port map( a => mult_125_ab_6_13_port, b => n1723, outb => n1722
                           );
   U1254 : nor2 port map( a => mult_125_ab_7_13_port, b => n1725, outb => n1724
                           );
   U1255 : nor2 port map( a => mult_125_ab_8_13_port, b => n1727, outb => n1726
                           );
   U1256 : nor2 port map( a => mult_125_ab_9_13_port, b => n1729, outb => n1728
                           );
   U1257 : nor2 port map( a => mult_125_ab_10_13_port, b => n1731, outb => 
                           n1730);
   U1258 : nor2 port map( a => mult_125_ab_11_13_port, b => n1733, outb => 
                           n1732);
   U1259 : nor2 port map( a => mult_125_ab_12_13_port, b => n1735, outb => 
                           n1734);
   U1260 : nor2 port map( a => mult_125_ab_13_13_port, b => n1737, outb => 
                           n1736);
   U1261 : nor2 port map( a => mult_125_ab_14_13_port, b => n1739, outb => 
                           n1738);
   U1262 : nor2 port map( a => mult_125_ab_15_13_port, b => n1741, outb => 
                           n1740);
   U1263 : nand2 port map( a => n1743, b => n1744, outb => n1742);
   U1264 : nor2 port map( a => mult_125_ab_3_12_port, b => n1746, outb => n1745
                           );
   U1265 : nor2 port map( a => mult_125_ab_4_12_port, b => n1748, outb => n1747
                           );
   U1266 : nor2 port map( a => mult_125_ab_5_12_port, b => n1750, outb => n1749
                           );
   U1267 : nor2 port map( a => mult_125_ab_6_12_port, b => n1752, outb => n1751
                           );
   U1268 : nor2 port map( a => mult_125_ab_7_12_port, b => n1754, outb => n1753
                           );
   U1269 : nor2 port map( a => mult_125_ab_8_12_port, b => n1756, outb => n1755
                           );
   U1270 : nor2 port map( a => mult_125_ab_9_12_port, b => n1758, outb => n1757
                           );
   U1271 : nor2 port map( a => mult_125_ab_10_12_port, b => n1760, outb => 
                           n1759);
   U1272 : nor2 port map( a => mult_125_ab_11_12_port, b => n1762, outb => 
                           n1761);
   U1273 : nor2 port map( a => mult_125_ab_12_12_port, b => n1764, outb => 
                           n1763);
   U1274 : nor2 port map( a => mult_125_ab_13_12_port, b => n1766, outb => 
                           n1765);
   U1275 : nor2 port map( a => mult_125_ab_14_12_port, b => n1768, outb => 
                           n1767);
   U1276 : nor2 port map( a => mult_125_ab_15_12_port, b => n1770, outb => 
                           n1769);
   U1277 : nand2 port map( a => n1772, b => n1773, outb => n1771);
   U1278 : nand2 port map( a => n1775, b => n1776, outb => n1774);
   U1279 : nor2 port map( a => mult_125_ab_4_11_port, b => n1778, outb => n1777
                           );
   U1280 : nor2 port map( a => mult_125_ab_5_11_port, b => n1780, outb => n1779
                           );
   U1281 : nor2 port map( a => mult_125_ab_6_11_port, b => n1782, outb => n1781
                           );
   U1282 : nor2 port map( a => mult_125_ab_7_11_port, b => n1784, outb => n1783
                           );
   U1283 : nor2 port map( a => mult_125_ab_8_11_port, b => n1786, outb => n1785
                           );
   U1284 : nor2 port map( a => mult_125_ab_9_11_port, b => n1788, outb => n1787
                           );
   U1285 : nor2 port map( a => mult_125_ab_10_11_port, b => n1790, outb => 
                           n1789);
   U1286 : nor2 port map( a => mult_125_ab_11_11_port, b => n1792, outb => 
                           n1791);
   U1287 : nor2 port map( a => mult_125_ab_12_11_port, b => n1794, outb => 
                           n1793);
   U1288 : nor2 port map( a => mult_125_ab_13_11_port, b => n1796, outb => 
                           n1795);
   U1289 : nor2 port map( a => mult_125_ab_14_11_port, b => n1798, outb => 
                           n1797);
   U1290 : nand2 port map( a => n1800, b => n1801, outb => n1799);
   U1291 : nand2 port map( a => n1803, b => n1804, outb => n1802);
   U1292 : nor2 port map( a => mult_125_ab_3_10_port, b => n1806, outb => n1805
                           );
   U1293 : nor2 port map( a => mult_125_ab_4_10_port, b => n1808, outb => n1807
                           );
   U1294 : nand2 port map( a => n1810, b => n1811, outb => n1809);
   U1295 : nor2 port map( a => mult_125_ab_6_10_port, b => n1813, outb => n1812
                           );
   U1296 : nor2 port map( a => mult_125_ab_7_10_port, b => n1815, outb => n1814
                           );
   U1297 : nor2 port map( a => mult_125_ab_8_10_port, b => n1817, outb => n1816
                           );
   U1298 : nor2 port map( a => mult_125_ab_9_10_port, b => n1819, outb => n1818
                           );
   U1299 : nor2 port map( a => mult_125_ab_10_10_port, b => n1821, outb => 
                           n1820);
   U1300 : nor2 port map( a => mult_125_ab_11_10_port, b => n1823, outb => 
                           n1822);
   U1301 : nor2 port map( a => mult_125_ab_12_10_port, b => n1825, outb => 
                           n1824);
   U1302 : nor2 port map( a => mult_125_ab_13_10_port, b => n1827, outb => 
                           n1826);
   U1303 : nor2 port map( a => mult_125_ab_14_10_port, b => n1829, outb => 
                           n1828);
   U1304 : nor2 port map( a => mult_125_ab_15_10_port, b => n1831, outb => 
                           n1830);
   U1305 : nand2 port map( a => n1833, b => n1834, outb => n1832);
   U1306 : nor2 port map( a => mult_125_ab_3_9_port, b => n1836, outb => n1835)
                           ;
   U1307 : nor2 port map( a => mult_125_ab_4_9_port, b => n1838, outb => n1837)
                           ;
   U1308 : nor2 port map( a => mult_125_ab_5_9_port, b => n1840, outb => n1839)
                           ;
   U1309 : nor2 port map( a => mult_125_ab_6_9_port, b => n1842, outb => n1841)
                           ;
   U1310 : nor2 port map( a => mult_125_ab_7_9_port, b => n1844, outb => n1843)
                           ;
   U1311 : nor2 port map( a => mult_125_ab_8_9_port, b => n1846, outb => n1845)
                           ;
   U1312 : nor2 port map( a => mult_125_ab_9_9_port, b => n1848, outb => n1847)
                           ;
   U1313 : nor2 port map( a => mult_125_ab_10_9_port, b => n1850, outb => n1849
                           );
   U1314 : nor2 port map( a => mult_125_ab_11_9_port, b => n1852, outb => n1851
                           );
   U1315 : nor2 port map( a => mult_125_ab_12_9_port, b => n1854, outb => n1853
                           );
   U1316 : nor2 port map( a => mult_125_ab_13_9_port, b => n1856, outb => n1855
                           );
   U1317 : nor2 port map( a => mult_125_ab_14_9_port, b => n1858, outb => n1857
                           );
   U1318 : nand2 port map( a => n1860, b => n1861, outb => n1859);
   U1319 : nand2 port map( a => n1863, b => n1864, outb => n1862);
   U1320 : nor2 port map( a => mult_125_ab_3_8_port, b => n1866, outb => n1865)
                           ;
   U1321 : nor2 port map( a => mult_125_ab_4_8_port, b => n1868, outb => n1867)
                           ;
   U1322 : nor2 port map( a => mult_125_ab_5_8_port, b => n1870, outb => n1869)
                           ;
   U1323 : nor2 port map( a => mult_125_ab_6_8_port, b => n1872, outb => n1871)
                           ;
   U1324 : nor2 port map( a => mult_125_ab_7_8_port, b => n1874, outb => n1873)
                           ;
   U1325 : nor2 port map( a => mult_125_ab_8_8_port, b => n1876, outb => n1875)
                           ;
   U1326 : nor2 port map( a => mult_125_ab_9_8_port, b => n1878, outb => n1877)
                           ;
   U1327 : nor2 port map( a => mult_125_ab_10_8_port, b => n1880, outb => n1879
                           );
   U1328 : nor2 port map( a => mult_125_ab_11_8_port, b => n1882, outb => n1881
                           );
   U1329 : nor2 port map( a => mult_125_ab_12_8_port, b => n1884, outb => n1883
                           );
   U1330 : nor2 port map( a => mult_125_ab_13_8_port, b => n1886, outb => n1885
                           );
   U1331 : nor2 port map( a => mult_125_ab_14_8_port, b => n1888, outb => n1887
                           );
   U1332 : nor2 port map( a => mult_125_ab_15_8_port, b => n1890, outb => n1889
                           );
   U1333 : nand2 port map( a => n1892, b => n1893, outb => n1891);
   U1334 : nand2 port map( a => n1895, b => n1896, outb => n1894);
   U1335 : nor2 port map( a => mult_125_ab_4_7_port, b => n1898, outb => n1897)
                           ;
   U1336 : nor2 port map( a => mult_125_ab_5_7_port, b => n1900, outb => n1899)
                           ;
   U1337 : nor2 port map( a => mult_125_ab_6_7_port, b => n1902, outb => n1901)
                           ;
   U1338 : nor2 port map( a => mult_125_ab_7_7_port, b => n1904, outb => n1903)
                           ;
   U1339 : nor2 port map( a => mult_125_ab_8_7_port, b => n1906, outb => n1905)
                           ;
   U1340 : nor2 port map( a => mult_125_ab_9_7_port, b => n1908, outb => n1907)
                           ;
   U1341 : nor2 port map( a => mult_125_ab_10_7_port, b => n1910, outb => n1909
                           );
   U1342 : nor2 port map( a => mult_125_ab_11_7_port, b => n1912, outb => n1911
                           );
   U1343 : nor2 port map( a => mult_125_ab_12_7_port, b => n1914, outb => n1913
                           );
   U1344 : nor2 port map( a => mult_125_ab_13_7_port, b => n1916, outb => n1915
                           );
   U1345 : nor2 port map( a => mult_125_ab_14_7_port, b => n1918, outb => n1917
                           );
   U1346 : nand2 port map( a => n1920, b => n1921, outb => n1919);
   U1347 : nand2 port map( a => n1923, b => n1924, outb => n1922);
   U1348 : nor2 port map( a => mult_125_ab_3_6_port, b => n1926, outb => n1925)
                           ;
   U1349 : nor2 port map( a => mult_125_ab_4_6_port, b => n1928, outb => n1927)
                           ;
   U1350 : nand2 port map( a => n1930, b => n1931, outb => n1929);
   U1351 : nor2 port map( a => mult_125_ab_6_6_port, b => n1933, outb => n1932)
                           ;
   U1352 : nor2 port map( a => mult_125_ab_7_6_port, b => n1935, outb => n1934)
                           ;
   U1353 : nor2 port map( a => mult_125_ab_8_6_port, b => n1937, outb => n1936)
                           ;
   U1354 : nand2 port map( a => n1939, b => n1940, outb => n1938);
   U1355 : nor2 port map( a => mult_125_ab_10_6_port, b => n1942, outb => n1941
                           );
   U1356 : nor2 port map( a => mult_125_ab_11_6_port, b => n1944, outb => n1943
                           );
   U1357 : nor2 port map( a => mult_125_ab_12_6_port, b => n1946, outb => n1945
                           );
   U1358 : nor2 port map( a => mult_125_ab_13_6_port, b => n1948, outb => n1947
                           );
   U1359 : nor2 port map( a => mult_125_ab_14_6_port, b => n1950, outb => n1949
                           );
   U1360 : nor2 port map( a => mult_125_ab_15_6_port, b => n1952, outb => n1951
                           );
   U1361 : nand2 port map( a => n1954, b => n1955, outb => n1953);
   U1362 : nand2 port map( a => n1957, b => n1958, outb => n1956);
   U1363 : nor2 port map( a => mult_125_ab_4_5_port, b => n1960, outb => n1959)
                           ;
   U1364 : nor2 port map( a => mult_125_ab_5_5_port, b => n1962, outb => n1961)
                           ;
   U1365 : nand2 port map( a => n1964, b => n1965, outb => n1963);
   U1366 : nor2 port map( a => mult_125_ab_7_5_port, b => n1967, outb => n1966)
                           ;
   U1367 : nor2 port map( a => mult_125_ab_8_5_port, b => n1969, outb => n1968)
                           ;
   U1368 : nor2 port map( a => mult_125_ab_9_5_port, b => n1971, outb => n1970)
                           ;
   U1369 : nor2 port map( a => mult_125_ab_10_5_port, b => n1973, outb => n1972
                           );
   U1370 : nor2 port map( a => mult_125_ab_11_5_port, b => n1975, outb => n1974
                           );
   U1371 : nor2 port map( a => mult_125_ab_12_5_port, b => n1977, outb => n1976
                           );
   U1372 : nor2 port map( a => mult_125_ab_13_5_port, b => n1979, outb => n1978
                           );
   U1373 : nor2 port map( a => mult_125_ab_14_5_port, b => n1981, outb => n1980
                           );
   U1374 : nand2 port map( a => n1983, b => n1984, outb => n1982);
   U1375 : nand2 port map( a => n1986, b => n1987, outb => n1985);
   U1376 : nor2 port map( a => mult_125_ab_3_4_port, b => n1989, outb => n1988)
                           ;
   U1377 : nor2 port map( a => mult_125_ab_4_4_port, b => n1991, outb => n1990)
                           ;
   U1378 : nand2 port map( a => n1993, b => n1994, outb => n1992);
   U1379 : nor2 port map( a => mult_125_ab_6_4_port, b => n1996, outb => n1995)
                           ;
   U1380 : nand2 port map( a => n1998, b => n1999, outb => n1997);
   U1381 : nor2 port map( a => mult_125_ab_8_4_port, b => n2001, outb => n2000)
                           ;
   U1382 : nor2 port map( a => mult_125_ab_9_4_port, b => n2003, outb => n2002)
                           ;
   U1383 : nor2 port map( a => mult_125_ab_10_4_port, b => n2005, outb => n2004
                           );
   U1384 : nand2 port map( a => n2007, b => n2008, outb => n2006);
   U1385 : nor2 port map( a => mult_125_ab_12_4_port, b => n2010, outb => n2009
                           );
   U1386 : nor2 port map( a => mult_125_ab_13_4_port, b => n2012, outb => n2011
                           );
   U1387 : nor2 port map( a => mult_125_ab_14_4_port, b => n2014, outb => n2013
                           );
   U1388 : nand2 port map( a => n2016, b => n2017, outb => n2015);
   U1389 : nand2 port map( a => n2019, b => n2020, outb => n2018);
   U1390 : nand2 port map( a => n2022, b => n2023, outb => n2021);
   U1391 : nor2 port map( a => mult_125_ab_4_3_port, b => n2025, outb => n2024)
                           ;
   U1392 : nor2 port map( a => mult_125_ab_5_3_port, b => n2027, outb => n2026)
                           ;
   U1393 : nor2 port map( a => mult_125_ab_6_3_port, b => n2029, outb => n2028)
                           ;
   U1394 : nor2 port map( a => mult_125_ab_7_3_port, b => n2031, outb => n2030)
                           ;
   U1395 : nor2 port map( a => mult_125_ab_8_3_port, b => n2033, outb => n2032)
                           ;
   U1396 : nor2 port map( a => mult_125_ab_9_3_port, b => n2035, outb => n2034)
                           ;
   U1397 : nor2 port map( a => mult_125_ab_10_3_port, b => n2037, outb => n2036
                           );
   U1398 : nor2 port map( a => mult_125_ab_11_3_port, b => n2039, outb => n2038
                           );
   U1399 : nor2 port map( a => mult_125_ab_12_3_port, b => n2041, outb => n2040
                           );
   U1400 : nor2 port map( a => mult_125_ab_13_3_port, b => n2043, outb => n2042
                           );
   U1401 : nor2 port map( a => mult_125_ab_14_3_port, b => n2045, outb => n2044
                           );
   U1402 : nor2 port map( a => mult_125_ab_15_3_port, b => n2047, outb => n2046
                           );
   U1403 : nand2 port map( a => n2049, b => n2050, outb => n2048);
   U1404 : nor2 port map( a => mult_125_ab_3_2_port, b => n2052, outb => n2051)
                           ;
   U1405 : nor2 port map( a => mult_125_ab_4_2_port, b => n2054, outb => n2053)
                           ;
   U1406 : nor2 port map( a => mult_125_ab_5_2_port, b => n2056, outb => n2055)
                           ;
   U1407 : nor2 port map( a => mult_125_ab_6_2_port, b => n2058, outb => n2057)
                           ;
   U1408 : nand2 port map( a => n2060, b => n2061, outb => n2059);
   U1409 : nor2 port map( a => mult_125_ab_8_2_port, b => n2063, outb => n2062)
                           ;
   U1410 : nor2 port map( a => mult_125_ab_9_2_port, b => n2065, outb => n2064)
                           ;
   U1411 : nor2 port map( a => mult_125_ab_10_2_port, b => n2067, outb => n2066
                           );
   U1412 : nor2 port map( a => mult_125_ab_11_2_port, b => n2069, outb => n2068
                           );
   U1413 : nor2 port map( a => mult_125_ab_12_2_port, b => n2071, outb => n2070
                           );
   U1414 : nor2 port map( a => mult_125_ab_13_2_port, b => n2073, outb => n2072
                           );
   U1415 : nor2 port map( a => mult_125_ab_14_2_port, b => n2075, outb => n2074
                           );
   U1416 : nor2 port map( a => mult_125_ab_15_2_port, b => n2077, outb => n2076
                           );
   U1417 : nand2 port map( a => n2079, b => n2080, outb => n2078);
   U1418 : nor2 port map( a => mult_125_ab_3_1_port, b => n2082, outb => n2081)
                           ;
   U1419 : nor2 port map( a => mult_125_ab_4_1_port, b => n2084, outb => n2083)
                           ;
   U1420 : nor2 port map( a => mult_125_ab_5_1_port, b => n2086, outb => n2085)
                           ;
   U1421 : nor2 port map( a => mult_125_ab_6_1_port, b => n2088, outb => n2087)
                           ;
   U1422 : nor2 port map( a => mult_125_ab_7_1_port, b => n2090, outb => n2089)
                           ;
   U1423 : nor2 port map( a => mult_125_ab_8_1_port, b => n2092, outb => n2091)
                           ;
   U1424 : nor2 port map( a => mult_125_ab_9_1_port, b => n2094, outb => n2093)
                           ;
   U1425 : nor2 port map( a => mult_125_ab_10_1_port, b => n2096, outb => n2095
                           );
   U1426 : nor2 port map( a => mult_125_ab_11_1_port, b => n2098, outb => n2097
                           );
   U1427 : nor2 port map( a => mult_125_ab_12_1_port, b => n2100, outb => n2099
                           );
   U1428 : nor2 port map( a => mult_125_ab_13_1_port, b => n2102, outb => n2101
                           );
   U1429 : nor2 port map( a => mult_125_ab_14_1_port, b => n2104, outb => n2103
                           );
   U1430 : nor2 port map( a => mult_125_ab_15_1_port, b => n2106, outb => n2105
                           );
   U1431 : nor2 port map( a => mult_125_ab_2_0_port, b => n2108, outb => n2107)
                           ;
   U1432 : nor2 port map( a => mult_125_ab_3_0_port, b => n2110, outb => n2109)
                           ;
   U1433 : nor2 port map( a => mult_125_ab_4_0_port, b => n2112, outb => n2111)
                           ;
   U1434 : nor2 port map( a => mult_125_ab_5_0_port, b => n2114, outb => n2113)
                           ;
   U1435 : nor2 port map( a => mult_125_ab_6_0_port, b => n2116, outb => n2115)
                           ;
   U1436 : nor2 port map( a => mult_125_ab_7_0_port, b => n2118, outb => n2117)
                           ;
   U1437 : nor2 port map( a => mult_125_ab_8_0_port, b => n2120, outb => n2119)
                           ;
   U1438 : nor2 port map( a => mult_125_ab_9_0_port, b => n2122, outb => n2121)
                           ;
   U1439 : nor2 port map( a => mult_125_ab_10_0_port, b => n2124, outb => n2123
                           );
   U1440 : nor2 port map( a => mult_125_ab_11_0_port, b => n2126, outb => n2125
                           );
   U1441 : nor2 port map( a => mult_125_ab_12_0_port, b => n2128, outb => n2127
                           );
   U1442 : nor2 port map( a => mult_125_ab_13_0_port, b => n2130, outb => n2129
                           );
   U1443 : nor2 port map( a => mult_125_ab_14_0_port, b => n2132, outb => n2131
                           );
   U1444 : nor2 port map( a => mult_125_ab_15_0_port, b => n2134, outb => n2133
                           );
   U1445 : nor2 port map( a => mult_125_ZB, b => mult_125_ZA, outb => n310);
   U1446 : nand2 port map( a => mult_125_QB, b => mult_125_ab_15_15_port, outb 
                           => n2135);
   U1447 : nor2 port map( a => adder_mem_array_3_1_port, b => n2137, outb => 
                           n2136);
   U1448 : nor2 port map( a => multiplier_sigs_2_2_port, b => 
                           adder_mem_array_3_2_port, outb => n2138);
   U1449 : nor2 port map( a => multiplier_sigs_2_3_port, b => 
                           adder_mem_array_3_3_port, outb => n2139);
   U1450 : nor2 port map( a => multiplier_sigs_2_4_port, b => 
                           adder_mem_array_3_4_port, outb => n2140);
   U1451 : nor2 port map( a => multiplier_sigs_2_5_port, b => 
                           adder_mem_array_3_5_port, outb => n2141);
   U1452 : nor2 port map( a => multiplier_sigs_2_6_port, b => 
                           adder_mem_array_3_6_port, outb => n2142);
   U1453 : nor2 port map( a => multiplier_sigs_2_7_port, b => 
                           adder_mem_array_3_7_port, outb => n2143);
   U1454 : nor2 port map( a => multiplier_sigs_2_8_port, b => 
                           adder_mem_array_3_8_port, outb => n2144);
   U1455 : nor2 port map( a => multiplier_sigs_2_9_port, b => 
                           adder_mem_array_3_9_port, outb => n2145);
   U1456 : nor2 port map( a => multiplier_sigs_2_10_port, b => 
                           adder_mem_array_3_10_port, outb => n2146);
   U1457 : nor2 port map( a => multiplier_sigs_2_11_port, b => 
                           adder_mem_array_3_11_port, outb => n2147);
   U1458 : nor2 port map( a => multiplier_sigs_2_12_port, b => 
                           adder_mem_array_3_12_port, outb => n2148);
   U1459 : nor2 port map( a => multiplier_sigs_2_13_port, b => 
                           adder_mem_array_3_13_port, outb => n2149);
   U1460 : nor2 port map( a => multiplier_sigs_2_14_port, b => 
                           adder_mem_array_3_14_port, outb => n2150);
   U1461 : nor2 port map( a => multiplier_sigs_2_15_port, b => 
                           adder_mem_array_3_15_port, outb => n2151);
   U1462 : nor2 port map( a => multiplier_sigs_2_16_port, b => 
                           adder_mem_array_3_16_port, outb => n2152);
   U1463 : nor2 port map( a => multiplier_sigs_2_17_port, b => 
                           adder_mem_array_3_17_port, outb => n2153);
   U1464 : nor2 port map( a => multiplier_sigs_2_18_port, b => 
                           adder_mem_array_3_18_port, outb => n2154);
   U1465 : nor2 port map( a => multiplier_sigs_2_19_port, b => 
                           adder_mem_array_3_19_port, outb => n2155);
   U1466 : nor2 port map( a => multiplier_sigs_2_20_port, b => 
                           adder_mem_array_3_20_port, outb => n2156);
   U1467 : nor2 port map( a => multiplier_sigs_2_21_port, b => 
                           adder_mem_array_3_21_port, outb => n2157);
   U1468 : nor2 port map( a => multiplier_sigs_2_22_port, b => 
                           adder_mem_array_3_22_port, outb => n2158);
   U1469 : nor2 port map( a => multiplier_sigs_2_23_port, b => 
                           adder_mem_array_3_23_port, outb => n2159);
   U1470 : nor2 port map( a => multiplier_sigs_2_24_port, b => 
                           adder_mem_array_3_24_port, outb => n2160);
   U1471 : nor2 port map( a => multiplier_sigs_2_25_port, b => 
                           adder_mem_array_3_25_port, outb => n2161);
   U1472 : nor2 port map( a => multiplier_sigs_2_26_port, b => 
                           adder_mem_array_3_26_port, outb => n2162);
   U1473 : nor2 port map( a => adder_mem_array_1_1_port, b => n2164, outb => 
                           n2163);
   U1474 : nor2 port map( a => multiplier_sigs_0_2_port, b => 
                           adder_mem_array_1_2_port, outb => n2165);
   U1475 : nor2 port map( a => adder_mem_array_2_1_port, b => n2167, outb => 
                           n2166);
   U1476 : nor2 port map( a => multiplier_sigs_1_2_port, b => 
                           adder_mem_array_2_2_port, outb => n2168);
   U1477 : nor2 port map( a => multiplier_sigs_1_3_port, b => 
                           adder_mem_array_2_3_port, outb => n2169);
   U1478 : nor2 port map( a => multiplier_sigs_1_4_port, b => 
                           adder_mem_array_2_4_port, outb => n2170);
   U1479 : nor2 port map( a => multiplier_sigs_1_5_port, b => 
                           adder_mem_array_2_5_port, outb => n2171);
   U1480 : nor2 port map( a => multiplier_sigs_1_6_port, b => 
                           adder_mem_array_2_6_port, outb => n2172);
   U1481 : nor2 port map( a => multiplier_sigs_1_7_port, b => 
                           adder_mem_array_2_7_port, outb => n2173);
   U1482 : nor2 port map( a => multiplier_sigs_1_8_port, b => 
                           adder_mem_array_2_8_port, outb => n2174);
   U1483 : nor2 port map( a => multiplier_sigs_1_9_port, b => 
                           adder_mem_array_2_9_port, outb => n2175);
   U1484 : nor2 port map( a => multiplier_sigs_1_10_port, b => 
                           adder_mem_array_2_10_port, outb => n2176);
   U1485 : nor2 port map( a => multiplier_sigs_1_11_port, b => 
                           adder_mem_array_2_11_port, outb => n2177);
   U1486 : nor2 port map( a => multiplier_sigs_1_12_port, b => 
                           adder_mem_array_2_12_port, outb => n2178);
   U1487 : nor2 port map( a => multiplier_sigs_1_13_port, b => 
                           adder_mem_array_2_13_port, outb => n2179);
   U1488 : nor2 port map( a => multiplier_sigs_1_14_port, b => 
                           adder_mem_array_2_14_port, outb => n2180);
   U1489 : nor2 port map( a => multiplier_sigs_1_15_port, b => 
                           adder_mem_array_2_15_port, outb => n2181);
   U1490 : nor2 port map( a => multiplier_sigs_1_16_port, b => 
                           adder_mem_array_2_16_port, outb => n2182);
   U1491 : nor2 port map( a => multiplier_sigs_1_17_port, b => 
                           adder_mem_array_2_17_port, outb => n2183);
   U1492 : nor2 port map( a => multiplier_sigs_1_18_port, b => 
                           adder_mem_array_2_18_port, outb => n2184);
   U1493 : nor2 port map( a => multiplier_sigs_1_19_port, b => 
                           adder_mem_array_2_19_port, outb => n2185);
   U1494 : nor2 port map( a => multiplier_sigs_1_20_port, b => 
                           adder_mem_array_2_20_port, outb => n2186);
   U1495 : nor2 port map( a => multiplier_sigs_1_21_port, b => 
                           adder_mem_array_2_21_port, outb => n2187);
   U1496 : nor2 port map( a => multiplier_sigs_1_22_port, b => 
                           adder_mem_array_2_22_port, outb => n2188);
   U1497 : nor2 port map( a => multiplier_sigs_1_23_port, b => 
                           adder_mem_array_2_23_port, outb => n2189);
   U1498 : nor2 port map( a => multiplier_sigs_1_24_port, b => 
                           adder_mem_array_2_24_port, outb => n2190);
   U1499 : nor2 port map( a => multiplier_sigs_1_25_port, b => 
                           adder_mem_array_2_25_port, outb => n2191);
   U1500 : nor2 port map( a => multiplier_sigs_1_26_port, b => 
                           adder_mem_array_2_26_port, outb => n2192);
   U1501 : nor2 port map( a => multiplier_sigs_1_27_port, b => 
                           adder_mem_array_2_27_port, outb => n2193);
   U1502 : nor2 port map( a => multiplier_sigs_1_28_port, b => 
                           adder_mem_array_2_28_port, outb => n2194);
   U1503 : nor2 port map( a => multiplier_sigs_1_29_port, b => 
                           adder_mem_array_2_29_port, outb => n2195);
   U1504 : nor2 port map( a => multiplier_sigs_1_30_port, b => 
                           adder_mem_array_2_30_port, outb => n2196);
   U1505 : aoi22 port map( a => n2198, b => n2199, c => 
                           adder_mem_array_2_31_port, d => 
                           multiplier_sigs_1_31_port, outb => n2197);
   U1506 : nor2 port map( a => multiplier_sigs_0_3_port, b => 
                           adder_mem_array_1_3_port, outb => n2200);
   U1507 : nor2 port map( a => multiplier_sigs_0_4_port, b => 
                           adder_mem_array_1_4_port, outb => n2201);
   U1508 : nor2 port map( a => multiplier_sigs_0_5_port, b => 
                           adder_mem_array_1_5_port, outb => n2202);
   U1509 : nor2 port map( a => multiplier_sigs_0_6_port, b => 
                           adder_mem_array_1_6_port, outb => n2203);
   U1510 : nor2 port map( a => multiplier_sigs_0_7_port, b => 
                           adder_mem_array_1_7_port, outb => n2204);
   U1511 : nor2 port map( a => multiplier_sigs_0_8_port, b => 
                           adder_mem_array_1_8_port, outb => n2205);
   U1512 : nor2 port map( a => multiplier_sigs_0_9_port, b => 
                           adder_mem_array_1_9_port, outb => n2206);
   U1513 : nor2 port map( a => multiplier_sigs_0_10_port, b => 
                           adder_mem_array_1_10_port, outb => n2207);
   U1514 : nor2 port map( a => multiplier_sigs_0_11_port, b => 
                           adder_mem_array_1_11_port, outb => n2208);
   U1515 : nor2 port map( a => multiplier_sigs_0_12_port, b => 
                           adder_mem_array_1_12_port, outb => n2209);
   U1516 : nor2 port map( a => multiplier_sigs_0_13_port, b => 
                           adder_mem_array_1_13_port, outb => n2210);
   U1517 : nor2 port map( a => multiplier_sigs_0_14_port, b => 
                           adder_mem_array_1_14_port, outb => n2211);
   U1518 : nor2 port map( a => multiplier_sigs_0_15_port, b => 
                           adder_mem_array_1_15_port, outb => n2212);
   U1519 : nor2 port map( a => multiplier_sigs_0_16_port, b => 
                           adder_mem_array_1_16_port, outb => n2213);
   U1520 : nor2 port map( a => multiplier_sigs_0_17_port, b => 
                           adder_mem_array_1_17_port, outb => n2214);
   U1521 : nor2 port map( a => multiplier_sigs_0_18_port, b => 
                           adder_mem_array_1_18_port, outb => n2215);
   U1522 : nor2 port map( a => multiplier_sigs_0_19_port, b => 
                           adder_mem_array_1_19_port, outb => n2216);
   U1523 : nor2 port map( a => multiplier_sigs_0_20_port, b => 
                           adder_mem_array_1_20_port, outb => n2217);
   U1524 : nor2 port map( a => multiplier_sigs_0_21_port, b => 
                           adder_mem_array_1_21_port, outb => n2218);
   U1525 : nor2 port map( a => multiplier_sigs_0_22_port, b => 
                           adder_mem_array_1_22_port, outb => n2219);
   U1526 : nor2 port map( a => multiplier_sigs_0_23_port, b => 
                           adder_mem_array_1_23_port, outb => n2220);
   U1527 : nor2 port map( a => multiplier_sigs_0_24_port, b => 
                           adder_mem_array_1_24_port, outb => n2221);
   U1528 : nor2 port map( a => multiplier_sigs_0_25_port, b => 
                           adder_mem_array_1_25_port, outb => n2222);
   U1529 : nor2 port map( a => multiplier_sigs_0_26_port, b => 
                           adder_mem_array_1_26_port, outb => n2223);
   U1530 : nor2 port map( a => multiplier_sigs_0_27_port, b => 
                           adder_mem_array_1_27_port, outb => n2224);
   U1531 : nor2 port map( a => multiplier_sigs_0_28_port, b => 
                           adder_mem_array_1_28_port, outb => n2225);
   U1532 : nor2 port map( a => multiplier_sigs_0_29_port, b => 
                           adder_mem_array_1_29_port, outb => n2226);
   U1533 : nor2 port map( a => multiplier_sigs_0_30_port, b => 
                           adder_mem_array_1_30_port, outb => n2227);
   U1534 : aoi22 port map( a => n2229, b => n2230, c => 
                           adder_mem_array_1_31_port, d => 
                           multiplier_sigs_0_31_port, outb => n2228);
   U1535 : nor2 port map( a => multiplier_sigs_2_27_port, b => 
                           adder_mem_array_3_27_port, outb => n2231);
   U1536 : nor2 port map( a => multiplier_sigs_2_28_port, b => 
                           adder_mem_array_3_28_port, outb => n2232);
   U1537 : nor2 port map( a => multiplier_sigs_2_29_port, b => 
                           adder_mem_array_3_29_port, outb => n2233);
   U1538 : nor2 port map( a => multiplier_sigs_2_30_port, b => 
                           adder_mem_array_3_30_port, outb => n2234);
   U1539 : aoi22 port map( a => n2236, b => n2237, c => 
                           adder_mem_array_3_31_port, d => 
                           multiplier_sigs_2_31_port, outb => n2235);
   U1540 : xor2 port map( a => mult_125_G4_ab_15_15_port, b => n2239, outb => 
                           n2238);
   U1541 : xor2 port map( a => mult_125_G4_ab_1_14_port, b => 
                           mult_125_G4_ab_0_15_port, outb => n2240);
   U1542 : xor2 port map( a => n2242, b => mult_125_G4_ab_1_15_port, outb => 
                           n2241);
   U1543 : xor2 port map( a => mult_125_G4_ab_1_13_port, b => 
                           mult_125_G4_ab_0_14_port, outb => n2243);
   U1544 : xor2 port map( a => n2245, b => n2240, outb => n2244);
   U1545 : xor2 port map( a => n2247, b => n2248, outb => n2246);
   U1546 : xor2 port map( a => n2250, b => n2251, outb => n2249);
   U1547 : xor2 port map( a => n2253, b => n2254, outb => n2252);
   U1548 : xor2 port map( a => n2256, b => n2257, outb => n2255);
   U1549 : xor2 port map( a => n2259, b => n2260, outb => n2258);
   U1550 : xor2 port map( a => n2262, b => n2263, outb => n2261);
   U1551 : xor2 port map( a => n2265, b => n2266, outb => n2264);
   U1552 : xor2 port map( a => n2268, b => n2269, outb => n2267);
   U1553 : xor2 port map( a => n2271, b => n2272, outb => n2270);
   U1554 : xor2 port map( a => n2274, b => n2275, outb => n2273);
   U1555 : xor2 port map( a => n2277, b => n2278, outb => n2276);
   U1556 : xor2 port map( a => n2279, b => n2280, outb => n246);
   U1557 : xor2 port map( a => mult_125_G4_ab_1_12_port, b => 
                           mult_125_G4_ab_0_13_port, outb => n2281);
   U1558 : xor2 port map( a => n2283, b => n2243, outb => n2282);
   U1559 : xor2 port map( a => n2285, b => n2286, outb => n2284);
   U1560 : xor2 port map( a => mult_125_G4_ab_1_11_port, b => 
                           mult_125_G4_ab_0_12_port, outb => n2287);
   U1561 : xor2 port map( a => n2289, b => n2281, outb => n2288);
   U1562 : xor2 port map( a => n2291, b => n2292, outb => n2290);
   U1563 : xor2 port map( a => n2294, b => n2295, outb => n2293);
   U1564 : xor2 port map( a => n2297, b => n2298, outb => n2296);
   U1565 : xor2 port map( a => n2300, b => n2301, outb => n2299);
   U1566 : xor2 port map( a => n2303, b => n2304, outb => n2302);
   U1567 : xor2 port map( a => n2306, b => n2307, outb => n2305);
   U1568 : xor2 port map( a => n2309, b => n2310, outb => n2308);
   U1569 : xor2 port map( a => n2312, b => n2313, outb => n2311);
   U1570 : xor2 port map( a => n2315, b => n2316, outb => n2314);
   U1571 : xor2 port map( a => n2318, b => n2319, outb => n2317);
   U1572 : xor2 port map( a => n2320, b => n2321, outb => n250);
   U1573 : xor2 port map( a => mult_125_G4_ab_1_10_port, b => 
                           mult_125_G4_ab_0_11_port, outb => n2322);
   U1574 : xor2 port map( a => n2324, b => n2287, outb => n2323);
   U1575 : xor2 port map( a => n2326, b => n2327, outb => n2325);
   U1576 : xor2 port map( a => n2329, b => n2330, outb => n2328);
   U1577 : xor2 port map( a => mult_125_G4_ab_1_9_port, b => 
                           mult_125_G4_ab_0_10_port, outb => n2331);
   U1578 : xor2 port map( a => n2333, b => n2322, outb => n2332);
   U1579 : xor2 port map( a => n2335, b => n2336, outb => n2334);
   U1580 : xor2 port map( a => n2338, b => n2339, outb => n2337);
   U1581 : xor2 port map( a => n2341, b => n2342, outb => n2340);
   U1582 : xor2 port map( a => n2344, b => n2345, outb => n2343);
   U1583 : xor2 port map( a => n2347, b => n2348, outb => n2346);
   U1584 : xor2 port map( a => n2350, b => n2351, outb => n2349);
   U1585 : xor2 port map( a => n2353, b => n2354, outb => n2352);
   U1586 : xor2 port map( a => n2356, b => n2357, outb => n2355);
   U1587 : xor2 port map( a => n2359, b => n2360, outb => n2358);
   U1588 : xor2 port map( a => n2361, b => n2362, outb => n254);
   U1589 : xor2 port map( a => mult_125_G4_ab_1_8_port, b => 
                           mult_125_G4_ab_0_9_port, outb => n2363);
   U1590 : xor2 port map( a => n2365, b => n2331, outb => n2364);
   U1591 : xor2 port map( a => n2367, b => n2368, outb => n2366);
   U1592 : xor2 port map( a => n2370, b => n2371, outb => n2369);
   U1593 : xor2 port map( a => n2373, b => n2374, outb => n2372);
   U1594 : xor2 port map( a => mult_125_G4_ab_1_7_port, b => 
                           mult_125_G4_ab_0_8_port, outb => n2375);
   U1595 : xor2 port map( a => n2377, b => n2363, outb => n2376);
   U1596 : xor2 port map( a => n2379, b => n2380, outb => n2378);
   U1597 : xor2 port map( a => n2382, b => n2383, outb => n2381);
   U1598 : xor2 port map( a => n2385, b => n2386, outb => n2384);
   U1599 : xor2 port map( a => n2388, b => n2389, outb => n2387);
   U1600 : xor2 port map( a => n2391, b => n2392, outb => n2390);
   U1601 : xor2 port map( a => n2394, b => n2395, outb => n2393);
   U1602 : xor2 port map( a => n2397, b => n2398, outb => n2396);
   U1603 : xor2 port map( a => n2400, b => n2401, outb => n2399);
   U1604 : xor2 port map( a => n2402, b => n2403, outb => n258);
   U1605 : xor2 port map( a => mult_125_G4_ab_1_6_port, b => 
                           mult_125_G4_ab_0_7_port, outb => n2404);
   U1606 : xor2 port map( a => n2406, b => n2375, outb => n2405);
   U1607 : xor2 port map( a => n2408, b => n2409, outb => n2407);
   U1608 : xor2 port map( a => n2411, b => n2412, outb => n2410);
   U1609 : xor2 port map( a => n2414, b => n2415, outb => n2413);
   U1610 : xor2 port map( a => n2417, b => n2418, outb => n2416);
   U1611 : xor2 port map( a => mult_125_G4_ab_1_5_port, b => 
                           mult_125_G4_ab_0_6_port, outb => n2419);
   U1612 : xor2 port map( a => n2421, b => n2404, outb => n2420);
   U1613 : xor2 port map( a => n2423, b => n2424, outb => n2422);
   U1614 : xor2 port map( a => n2426, b => n2427, outb => n2425);
   U1615 : xor2 port map( a => n2429, b => n2430, outb => n2428);
   U1616 : xor2 port map( a => n2432, b => n2433, outb => n2431);
   U1617 : xor2 port map( a => n2435, b => n2436, outb => n2434);
   U1618 : xor2 port map( a => n2438, b => n2439, outb => n2437);
   U1619 : xor2 port map( a => n2441, b => n2442, outb => n2440);
   U1620 : xor2 port map( a => n2443, b => n2444, outb => n262);
   U1621 : xor2 port map( a => mult_125_G4_ab_1_4_port, b => 
                           mult_125_G4_ab_0_5_port, outb => n2445);
   U1622 : xor2 port map( a => n2447, b => n2419, outb => n2446);
   U1623 : xor2 port map( a => n2449, b => n2450, outb => n2448);
   U1624 : xor2 port map( a => n2452, b => n2453, outb => n2451);
   U1625 : xor2 port map( a => n2455, b => n2456, outb => n2454);
   U1626 : xor2 port map( a => n2458, b => n2459, outb => n2457);
   U1627 : xor2 port map( a => n2461, b => n2462, outb => n2460);
   U1628 : xor2 port map( a => mult_125_G4_ab_1_3_port, b => 
                           mult_125_G4_ab_0_4_port, outb => n2463);
   U1629 : xor2 port map( a => n2465, b => n2445, outb => n2464);
   U1630 : xor2 port map( a => n2467, b => n2468, outb => n2466);
   U1631 : xor2 port map( a => n2470, b => n2471, outb => n2469);
   U1632 : xor2 port map( a => n2473, b => n2474, outb => n2472);
   U1633 : xor2 port map( a => n2476, b => n2477, outb => n2475);
   U1634 : xor2 port map( a => n2479, b => n2480, outb => n2478);
   U1635 : xor2 port map( a => n2482, b => n2483, outb => n2481);
   U1636 : xor2 port map( a => n2484, b => n2485, outb => n267);
   U1637 : xor2 port map( a => mult_125_G4_ab_1_2_port, b => 
                           mult_125_G4_ab_0_3_port, outb => n2486);
   U1638 : xor2 port map( a => n2488, b => n2463, outb => n2487);
   U1639 : xor2 port map( a => n2490, b => n2491, outb => n2489);
   U1640 : xor2 port map( a => n2493, b => n2494, outb => n2492);
   U1641 : xor2 port map( a => n2496, b => n2497, outb => n2495);
   U1642 : xor2 port map( a => n2499, b => n2500, outb => n2498);
   U1643 : xor2 port map( a => n2502, b => n2503, outb => n2501);
   U1644 : xor2 port map( a => n2505, b => n2506, outb => n2504);
   U1645 : xor2 port map( a => mult_125_G4_ab_1_1_port, b => 
                           mult_125_G4_ab_0_2_port, outb => n2507);
   U1646 : xor2 port map( a => n2509, b => n2486, outb => n2508);
   U1647 : xor2 port map( a => n2511, b => n2512, outb => n2510);
   U1648 : xor2 port map( a => n2514, b => n2515, outb => n2513);
   U1649 : xor2 port map( a => n2517, b => n2518, outb => n2516);
   U1650 : xor2 port map( a => n2520, b => n2521, outb => n2519);
   U1651 : xor2 port map( a => n2523, b => n2524, outb => n2522);
   U1652 : xor2 port map( a => n2526, b => n2527, outb => n2525);
   U1653 : xor2 port map( a => n2528, b => n2519, outb => mult_125_G4_A1_9_port
                           );
   U1654 : xor2 port map( a => n2529, b => n2516, outb => mult_125_G4_A1_7_port
                           );
   U1655 : xor2 port map( a => n2530, b => n2513, outb => mult_125_G4_A1_5_port
                           );
   U1656 : xor2 port map( a => n2531, b => n2510, outb => mult_125_G4_A1_3_port
                           );
   U1657 : xor2 port map( a => n242, b => n241, outb => mult_125_G4_A1_28_port)
                           ;
   U1658 : xor2 port map( a => n246, b => n245, outb => mult_125_G4_A1_26_port)
                           ;
   U1659 : xor2 port map( a => n250, b => n249, outb => mult_125_G4_A1_24_port)
                           ;
   U1660 : xor2 port map( a => n254, b => n253, outb => mult_125_G4_A1_22_port)
                           ;
   U1661 : xor2 port map( a => n258, b => n257, outb => mult_125_G4_A1_20_port)
                           ;
   U1662 : xor2 port map( a => n2532, b => n2508, outb => mult_125_G4_A1_1_port
                           );
   U1663 : xor2 port map( a => n262, b => n261, outb => mult_125_G4_A1_18_port)
                           ;
   U1664 : xor2 port map( a => n267, b => n266, outb => mult_125_G4_A1_16_port)
                           ;
   U1665 : xor2 port map( a => n2533, b => n275, outb => mult_125_G4_A1_13_port
                           );
   U1666 : xor2 port map( a => n2534, b => n2522, outb => 
                           mult_125_G4_A1_11_port);
   U1667 : xor2 port map( a => mult_125_G3_ab_15_15_port, b => n2536, outb => 
                           n2535);
   U1668 : xor2 port map( a => mult_125_G3_ab_1_14_port, b => 
                           mult_125_G3_ab_0_15_port, outb => n2537);
   U1669 : xor2 port map( a => n2539, b => mult_125_G3_ab_1_15_port, outb => 
                           n2538);
   U1670 : xor2 port map( a => mult_125_G3_ab_1_13_port, b => 
                           mult_125_G3_ab_0_14_port, outb => n2540);
   U1671 : xor2 port map( a => n2542, b => n2537, outb => n2541);
   U1672 : xor2 port map( a => n2544, b => n2545, outb => n2543);
   U1673 : xor2 port map( a => n2547, b => n2548, outb => n2546);
   U1674 : xor2 port map( a => n2550, b => n2551, outb => n2549);
   U1675 : xor2 port map( a => n2553, b => n2554, outb => n2552);
   U1676 : xor2 port map( a => n2556, b => n2557, outb => n2555);
   U1677 : xor2 port map( a => n2559, b => n2560, outb => n2558);
   U1678 : xor2 port map( a => n2562, b => n2563, outb => n2561);
   U1679 : xor2 port map( a => n2565, b => n2566, outb => n2564);
   U1680 : xor2 port map( a => n2568, b => n2569, outb => n2567);
   U1681 : xor2 port map( a => n2571, b => n2572, outb => n2570);
   U1682 : xor2 port map( a => n2574, b => n2575, outb => n2573);
   U1683 : xor2 port map( a => n2576, b => n2577, outb => n354);
   U1684 : xor2 port map( a => mult_125_G3_ab_1_12_port, b => 
                           mult_125_G3_ab_0_13_port, outb => n2578);
   U1685 : xor2 port map( a => n2580, b => n2540, outb => n2579);
   U1686 : xor2 port map( a => n2582, b => n2583, outb => n2581);
   U1687 : xor2 port map( a => mult_125_G3_ab_1_11_port, b => 
                           mult_125_G3_ab_0_12_port, outb => n2584);
   U1688 : xor2 port map( a => n2586, b => n2578, outb => n2585);
   U1689 : xor2 port map( a => n2588, b => n2589, outb => n2587);
   U1690 : xor2 port map( a => n2591, b => n2592, outb => n2590);
   U1691 : xor2 port map( a => n2594, b => n2595, outb => n2593);
   U1692 : xor2 port map( a => n2597, b => n2598, outb => n2596);
   U1693 : xor2 port map( a => n2600, b => n2601, outb => n2599);
   U1694 : xor2 port map( a => n2603, b => n2604, outb => n2602);
   U1695 : xor2 port map( a => n2606, b => n2607, outb => n2605);
   U1696 : xor2 port map( a => n2609, b => n2610, outb => n2608);
   U1697 : xor2 port map( a => n2612, b => n2613, outb => n2611);
   U1698 : xor2 port map( a => n2615, b => n2616, outb => n2614);
   U1699 : xor2 port map( a => n2617, b => n2618, outb => n358);
   U1700 : xor2 port map( a => mult_125_G3_ab_1_10_port, b => 
                           mult_125_G3_ab_0_11_port, outb => n2619);
   U1701 : xor2 port map( a => n2621, b => n2584, outb => n2620);
   U1702 : xor2 port map( a => n2623, b => n2624, outb => n2622);
   U1703 : xor2 port map( a => n2626, b => n2627, outb => n2625);
   U1704 : xor2 port map( a => mult_125_G3_ab_1_9_port, b => 
                           mult_125_G3_ab_0_10_port, outb => n2628);
   U1705 : xor2 port map( a => n2630, b => n2619, outb => n2629);
   U1706 : xor2 port map( a => n2632, b => n2633, outb => n2631);
   U1707 : xor2 port map( a => n2635, b => n2636, outb => n2634);
   U1708 : xor2 port map( a => n2638, b => n2639, outb => n2637);
   U1709 : xor2 port map( a => n2641, b => n2642, outb => n2640);
   U1710 : xor2 port map( a => n2644, b => n2645, outb => n2643);
   U1711 : xor2 port map( a => n2647, b => n2648, outb => n2646);
   U1712 : xor2 port map( a => n2650, b => n2651, outb => n2649);
   U1713 : xor2 port map( a => n2653, b => n2654, outb => n2652);
   U1714 : xor2 port map( a => n2656, b => n2657, outb => n2655);
   U1715 : xor2 port map( a => n2658, b => n2659, outb => n362);
   U1716 : xor2 port map( a => mult_125_G3_ab_1_8_port, b => 
                           mult_125_G3_ab_0_9_port, outb => n2660);
   U1717 : xor2 port map( a => n2662, b => n2628, outb => n2661);
   U1718 : xor2 port map( a => n2664, b => n2665, outb => n2663);
   U1719 : xor2 port map( a => n2667, b => n2668, outb => n2666);
   U1720 : xor2 port map( a => n2670, b => n2671, outb => n2669);
   U1721 : xor2 port map( a => mult_125_G3_ab_1_7_port, b => 
                           mult_125_G3_ab_0_8_port, outb => n2672);
   U1722 : xor2 port map( a => n2674, b => n2660, outb => n2673);
   U1723 : xor2 port map( a => n2676, b => n2677, outb => n2675);
   U1724 : xor2 port map( a => n2679, b => n2680, outb => n2678);
   U1725 : xor2 port map( a => n2682, b => n2683, outb => n2681);
   U1726 : xor2 port map( a => n2685, b => n2686, outb => n2684);
   U1727 : xor2 port map( a => n2688, b => n2689, outb => n2687);
   U1728 : xor2 port map( a => n2691, b => n2692, outb => n2690);
   U1729 : xor2 port map( a => n2694, b => n2695, outb => n2693);
   U1730 : xor2 port map( a => n2697, b => n2698, outb => n2696);
   U1731 : xor2 port map( a => n2699, b => n2700, outb => n366);
   U1732 : xor2 port map( a => mult_125_G3_ab_1_6_port, b => 
                           mult_125_G3_ab_0_7_port, outb => n2701);
   U1733 : xor2 port map( a => n2703, b => n2672, outb => n2702);
   U1734 : xor2 port map( a => n2705, b => n2706, outb => n2704);
   U1735 : xor2 port map( a => n2708, b => n2709, outb => n2707);
   U1736 : xor2 port map( a => n2711, b => n2712, outb => n2710);
   U1737 : xor2 port map( a => n2714, b => n2715, outb => n2713);
   U1738 : xor2 port map( a => mult_125_G3_ab_1_5_port, b => 
                           mult_125_G3_ab_0_6_port, outb => n2716);
   U1739 : xor2 port map( a => n2718, b => n2701, outb => n2717);
   U1740 : xor2 port map( a => n2720, b => n2721, outb => n2719);
   U1741 : xor2 port map( a => n2723, b => n2724, outb => n2722);
   U1742 : xor2 port map( a => n2726, b => n2727, outb => n2725);
   U1743 : xor2 port map( a => n2729, b => n2730, outb => n2728);
   U1744 : xor2 port map( a => n2732, b => n2733, outb => n2731);
   U1745 : xor2 port map( a => n2735, b => n2736, outb => n2734);
   U1746 : xor2 port map( a => n2738, b => n2739, outb => n2737);
   U1747 : xor2 port map( a => n2740, b => n2741, outb => n370);
   U1748 : xor2 port map( a => mult_125_G3_ab_1_4_port, b => 
                           mult_125_G3_ab_0_5_port, outb => n2742);
   U1749 : xor2 port map( a => n2744, b => n2716, outb => n2743);
   U1750 : xor2 port map( a => n2746, b => n2747, outb => n2745);
   U1751 : xor2 port map( a => n2749, b => n2750, outb => n2748);
   U1752 : xor2 port map( a => n2752, b => n2753, outb => n2751);
   U1753 : xor2 port map( a => n2755, b => n2756, outb => n2754);
   U1754 : xor2 port map( a => n2758, b => n2759, outb => n2757);
   U1755 : xor2 port map( a => mult_125_G3_ab_1_3_port, b => 
                           mult_125_G3_ab_0_4_port, outb => n2760);
   U1756 : xor2 port map( a => n2762, b => n2742, outb => n2761);
   U1757 : xor2 port map( a => n2764, b => n2765, outb => n2763);
   U1758 : xor2 port map( a => n2767, b => n2768, outb => n2766);
   U1759 : xor2 port map( a => n2770, b => n2771, outb => n2769);
   U1760 : xor2 port map( a => n2773, b => n2774, outb => n2772);
   U1761 : xor2 port map( a => n2776, b => n2777, outb => n2775);
   U1762 : xor2 port map( a => n2779, b => n2780, outb => n2778);
   U1763 : xor2 port map( a => n2781, b => n2782, outb => n375);
   U1764 : xor2 port map( a => mult_125_G3_ab_1_2_port, b => 
                           mult_125_G3_ab_0_3_port, outb => n2783);
   U1765 : xor2 port map( a => n2785, b => n2760, outb => n2784);
   U1766 : xor2 port map( a => n2787, b => n2788, outb => n2786);
   U1767 : xor2 port map( a => n2790, b => n2791, outb => n2789);
   U1768 : xor2 port map( a => n2793, b => n2794, outb => n2792);
   U1769 : xor2 port map( a => n2796, b => n2797, outb => n2795);
   U1770 : xor2 port map( a => n2799, b => n2800, outb => n2798);
   U1771 : xor2 port map( a => n2802, b => n2803, outb => n2801);
   U1772 : xor2 port map( a => mult_125_G3_ab_1_1_port, b => 
                           mult_125_G3_ab_0_2_port, outb => n2804);
   U1773 : xor2 port map( a => n2806, b => n2783, outb => n2805);
   U1774 : xor2 port map( a => n2808, b => n2809, outb => n2807);
   U1775 : xor2 port map( a => n2811, b => n2812, outb => n2810);
   U1776 : xor2 port map( a => n2814, b => n2815, outb => n2813);
   U1777 : xor2 port map( a => n2817, b => n2818, outb => n2816);
   U1778 : xor2 port map( a => n2820, b => n2821, outb => n2819);
   U1779 : xor2 port map( a => n2823, b => n2824, outb => n2822);
   U1780 : xor2 port map( a => n2825, b => n2816, outb => mult_125_G3_A1_9_port
                           );
   U1781 : xor2 port map( a => n2826, b => n2813, outb => mult_125_G3_A1_7_port
                           );
   U1782 : xor2 port map( a => n2827, b => n2810, outb => mult_125_G3_A1_5_port
                           );
   U1783 : xor2 port map( a => n2828, b => n2807, outb => mult_125_G3_A1_3_port
                           );
   U1784 : xor2 port map( a => n350, b => n349, outb => mult_125_G3_A1_28_port)
                           ;
   U1785 : xor2 port map( a => n354, b => n353, outb => mult_125_G3_A1_26_port)
                           ;
   U1786 : xor2 port map( a => n358, b => n357, outb => mult_125_G3_A1_24_port)
                           ;
   U1787 : xor2 port map( a => n362, b => n361, outb => mult_125_G3_A1_22_port)
                           ;
   U1788 : xor2 port map( a => n366, b => n365, outb => mult_125_G3_A1_20_port)
                           ;
   U1789 : xor2 port map( a => n2829, b => n2805, outb => mult_125_G3_A1_1_port
                           );
   U1790 : xor2 port map( a => n370, b => n369, outb => mult_125_G3_A1_18_port)
                           ;
   U1791 : xor2 port map( a => n375, b => n374, outb => mult_125_G3_A1_16_port)
                           ;
   U1792 : xor2 port map( a => n2830, b => n383, outb => mult_125_G3_A1_13_port
                           );
   U1793 : xor2 port map( a => n2831, b => n2819, outb => 
                           mult_125_G3_A1_11_port);
   U1794 : xor2 port map( a => mult_125_G2_ab_15_15_port, b => n2833, outb => 
                           n2832);
   U1795 : xor2 port map( a => mult_125_G2_ab_1_14_port, b => 
                           mult_125_G2_ab_0_15_port, outb => n2834);
   U1796 : xor2 port map( a => n2836, b => mult_125_G2_ab_1_15_port, outb => 
                           n2835);
   U1797 : xor2 port map( a => mult_125_G2_ab_1_13_port, b => 
                           mult_125_G2_ab_0_14_port, outb => n2837);
   U1798 : xor2 port map( a => n2839, b => n2834, outb => n2838);
   U1799 : xor2 port map( a => n2841, b => n2842, outb => n2840);
   U1800 : xor2 port map( a => n2844, b => n2845, outb => n2843);
   U1801 : xor2 port map( a => n2847, b => n2848, outb => n2846);
   U1802 : xor2 port map( a => n2850, b => n2851, outb => n2849);
   U1803 : xor2 port map( a => n2853, b => n2854, outb => n2852);
   U1804 : xor2 port map( a => n2856, b => n2857, outb => n2855);
   U1805 : xor2 port map( a => n2859, b => n2860, outb => n2858);
   U1806 : xor2 port map( a => n2862, b => n2863, outb => n2861);
   U1807 : xor2 port map( a => n2865, b => n2866, outb => n2864);
   U1808 : xor2 port map( a => n2868, b => n2869, outb => n2867);
   U1809 : xor2 port map( a => n2871, b => n2872, outb => n2870);
   U1810 : xor2 port map( a => n2873, b => n2874, outb => n318);
   U1811 : xor2 port map( a => mult_125_G2_ab_1_12_port, b => 
                           mult_125_G2_ab_0_13_port, outb => n2875);
   U1812 : xor2 port map( a => n2877, b => n2837, outb => n2876);
   U1813 : xor2 port map( a => n2879, b => n2880, outb => n2878);
   U1814 : xor2 port map( a => mult_125_G2_ab_1_11_port, b => 
                           mult_125_G2_ab_0_12_port, outb => n2881);
   U1815 : xor2 port map( a => n2883, b => n2875, outb => n2882);
   U1816 : xor2 port map( a => n2885, b => n2886, outb => n2884);
   U1817 : xor2 port map( a => n2888, b => n2889, outb => n2887);
   U1818 : xor2 port map( a => n2891, b => n2892, outb => n2890);
   U1819 : xor2 port map( a => n2894, b => n2895, outb => n2893);
   U1820 : xor2 port map( a => n2897, b => n2898, outb => n2896);
   U1821 : xor2 port map( a => n2900, b => n2901, outb => n2899);
   U1822 : xor2 port map( a => n2903, b => n2904, outb => n2902);
   U1823 : xor2 port map( a => n2906, b => n2907, outb => n2905);
   U1824 : xor2 port map( a => n2909, b => n2910, outb => n2908);
   U1825 : xor2 port map( a => n2912, b => n2913, outb => n2911);
   U1826 : xor2 port map( a => n2914, b => n2915, outb => n322);
   U1827 : xor2 port map( a => mult_125_G2_ab_1_10_port, b => 
                           mult_125_G2_ab_0_11_port, outb => n2916);
   U1828 : xor2 port map( a => n2918, b => n2881, outb => n2917);
   U1829 : xor2 port map( a => n2920, b => n2921, outb => n2919);
   U1830 : xor2 port map( a => n2923, b => n2924, outb => n2922);
   U1831 : xor2 port map( a => mult_125_G2_ab_1_9_port, b => 
                           mult_125_G2_ab_0_10_port, outb => n2925);
   U1832 : xor2 port map( a => n2927, b => n2916, outb => n2926);
   U1833 : xor2 port map( a => n2929, b => n2930, outb => n2928);
   U1834 : xor2 port map( a => n2932, b => n2933, outb => n2931);
   U1835 : xor2 port map( a => n2935, b => n2936, outb => n2934);
   U1836 : xor2 port map( a => n2938, b => n2939, outb => n2937);
   U1837 : xor2 port map( a => n2941, b => n2942, outb => n2940);
   U1838 : xor2 port map( a => n2944, b => n2945, outb => n2943);
   U1839 : xor2 port map( a => n2947, b => n2948, outb => n2946);
   U1840 : xor2 port map( a => n2950, b => n2951, outb => n2949);
   U1841 : xor2 port map( a => n2953, b => n2954, outb => n2952);
   U1842 : xor2 port map( a => n2955, b => n2956, outb => n326);
   U1843 : xor2 port map( a => mult_125_G2_ab_1_8_port, b => 
                           mult_125_G2_ab_0_9_port, outb => n2957);
   U1844 : xor2 port map( a => n2959, b => n2925, outb => n2958);
   U1845 : xor2 port map( a => n2961, b => n2962, outb => n2960);
   U1846 : xor2 port map( a => n2964, b => n2965, outb => n2963);
   U1847 : xor2 port map( a => n2967, b => n2968, outb => n2966);
   U1848 : xor2 port map( a => mult_125_G2_ab_1_7_port, b => 
                           mult_125_G2_ab_0_8_port, outb => n2969);
   U1849 : xor2 port map( a => n2971, b => n2957, outb => n2970);
   U1850 : xor2 port map( a => n2973, b => n2974, outb => n2972);
   U1851 : xor2 port map( a => n2976, b => n2977, outb => n2975);
   U1852 : xor2 port map( a => n2979, b => n2980, outb => n2978);
   U1853 : xor2 port map( a => n2982, b => n2983, outb => n2981);
   U1854 : xor2 port map( a => n2985, b => n2986, outb => n2984);
   U1855 : xor2 port map( a => n2988, b => n2989, outb => n2987);
   U1856 : xor2 port map( a => n2991, b => n2992, outb => n2990);
   U1857 : xor2 port map( a => n2994, b => n2995, outb => n2993);
   U1858 : xor2 port map( a => n2996, b => n2997, outb => n330);
   U1859 : xor2 port map( a => mult_125_G2_ab_1_6_port, b => 
                           mult_125_G2_ab_0_7_port, outb => n2998);
   U1860 : xor2 port map( a => n3000, b => n2969, outb => n2999);
   U1861 : xor2 port map( a => n3002, b => n3003, outb => n3001);
   U1862 : xor2 port map( a => n3005, b => n3006, outb => n3004);
   U1863 : xor2 port map( a => n3008, b => n3009, outb => n3007);
   U1864 : xor2 port map( a => n3011, b => n3012, outb => n3010);
   U1865 : xor2 port map( a => mult_125_G2_ab_1_5_port, b => 
                           mult_125_G2_ab_0_6_port, outb => n3013);
   U1866 : xor2 port map( a => n3015, b => n2998, outb => n3014);
   U1867 : xor2 port map( a => n3017, b => n3018, outb => n3016);
   U1868 : xor2 port map( a => n3020, b => n3021, outb => n3019);
   U1869 : xor2 port map( a => n3023, b => n3024, outb => n3022);
   U1870 : xor2 port map( a => n3026, b => n3027, outb => n3025);
   U1871 : xor2 port map( a => n3029, b => n3030, outb => n3028);
   U1872 : xor2 port map( a => n3032, b => n3033, outb => n3031);
   U1873 : xor2 port map( a => n3035, b => n3036, outb => n3034);
   U1874 : xor2 port map( a => n3037, b => n3038, outb => n334);
   U1875 : xor2 port map( a => mult_125_G2_ab_1_4_port, b => 
                           mult_125_G2_ab_0_5_port, outb => n3039);
   U1876 : xor2 port map( a => n3041, b => n3013, outb => n3040);
   U1877 : xor2 port map( a => n3043, b => n3044, outb => n3042);
   U1878 : xor2 port map( a => n3046, b => n3047, outb => n3045);
   U1879 : xor2 port map( a => n3049, b => n3050, outb => n3048);
   U1880 : xor2 port map( a => n3052, b => n3053, outb => n3051);
   U1881 : xor2 port map( a => n3055, b => n3056, outb => n3054);
   U1882 : xor2 port map( a => mult_125_G2_ab_1_3_port, b => 
                           mult_125_G2_ab_0_4_port, outb => n3057);
   U1883 : xor2 port map( a => n3059, b => n3039, outb => n3058);
   U1884 : xor2 port map( a => n3061, b => n3062, outb => n3060);
   U1885 : xor2 port map( a => n3064, b => n3065, outb => n3063);
   U1886 : xor2 port map( a => n3067, b => n3068, outb => n3066);
   U1887 : xor2 port map( a => n3070, b => n3071, outb => n3069);
   U1888 : xor2 port map( a => n3073, b => n3074, outb => n3072);
   U1889 : xor2 port map( a => n3076, b => n3077, outb => n3075);
   U1890 : xor2 port map( a => n3078, b => n3079, outb => n339);
   U1891 : xor2 port map( a => mult_125_G2_ab_1_2_port, b => 
                           mult_125_G2_ab_0_3_port, outb => n3080);
   U1892 : xor2 port map( a => n3082, b => n3057, outb => n3081);
   U1893 : xor2 port map( a => n3084, b => n3085, outb => n3083);
   U1894 : xor2 port map( a => n3087, b => n3088, outb => n3086);
   U1895 : xor2 port map( a => n3090, b => n3091, outb => n3089);
   U1896 : xor2 port map( a => n3093, b => n3094, outb => n3092);
   U1897 : xor2 port map( a => n3096, b => n3097, outb => n3095);
   U1898 : xor2 port map( a => n3099, b => n3100, outb => n3098);
   U1899 : xor2 port map( a => mult_125_G2_ab_1_1_port, b => 
                           mult_125_G2_ab_0_2_port, outb => n3101);
   U1900 : xor2 port map( a => n3103, b => n3080, outb => n3102);
   U1901 : xor2 port map( a => n3105, b => n3106, outb => n3104);
   U1902 : xor2 port map( a => n3108, b => n3109, outb => n3107);
   U1903 : xor2 port map( a => n3111, b => n3112, outb => n3110);
   U1904 : xor2 port map( a => n3114, b => n3115, outb => n3113);
   U1905 : xor2 port map( a => n3117, b => n3118, outb => n3116);
   U1906 : xor2 port map( a => n3120, b => n3121, outb => n3119);
   U1907 : xor2 port map( a => n3122, b => n3113, outb => mult_125_G2_A1_9_port
                           );
   U1908 : xor2 port map( a => n3123, b => n3110, outb => mult_125_G2_A1_7_port
                           );
   U1909 : xor2 port map( a => n3124, b => n3107, outb => mult_125_G2_A1_5_port
                           );
   U1910 : xor2 port map( a => n3125, b => n3104, outb => mult_125_G2_A1_3_port
                           );
   U1911 : xor2 port map( a => n314, b => n313, outb => mult_125_G2_A1_28_port)
                           ;
   U1912 : xor2 port map( a => n318, b => n317, outb => mult_125_G2_A1_26_port)
                           ;
   U1913 : xor2 port map( a => n322, b => n321, outb => mult_125_G2_A1_24_port)
                           ;
   U1914 : xor2 port map( a => n326, b => n325, outb => mult_125_G2_A1_22_port)
                           ;
   U1915 : xor2 port map( a => n330, b => n329, outb => mult_125_G2_A1_20_port)
                           ;
   U1916 : xor2 port map( a => n3126, b => n3102, outb => mult_125_G2_A1_1_port
                           );
   U1917 : xor2 port map( a => n334, b => n333, outb => mult_125_G2_A1_18_port)
                           ;
   U1918 : xor2 port map( a => n339, b => n338, outb => mult_125_G2_A1_16_port)
                           ;
   U1919 : xor2 port map( a => n3127, b => n347, outb => mult_125_G2_A1_13_port
                           );
   U1920 : xor2 port map( a => n3128, b => n3116, outb => 
                           mult_125_G2_A1_11_port);
   U1921 : xor2 port map( a => mult_125_ab_15_15_port, b => n3130, outb => 
                           n3129);
   U1922 : xor2 port map( a => mult_125_ab_1_14_port, b => 
                           mult_125_ab_0_15_port, outb => n3131);
   U1923 : xor2 port map( a => n3133, b => mult_125_ab_1_15_port, outb => n3132
                           );
   U1924 : xor2 port map( a => mult_125_ab_1_13_port, b => 
                           mult_125_ab_0_14_port, outb => n3134);
   U1925 : xor2 port map( a => n3136, b => n3131, outb => n3135);
   U1926 : xor2 port map( a => n3138, b => n3139, outb => n3137);
   U1927 : xor2 port map( a => n3141, b => n3142, outb => n3140);
   U1928 : xor2 port map( a => n3144, b => n3145, outb => n3143);
   U1929 : xor2 port map( a => n3147, b => n3148, outb => n3146);
   U1930 : xor2 port map( a => n3150, b => n3151, outb => n3149);
   U1931 : xor2 port map( a => n3153, b => n3154, outb => n3152);
   U1932 : xor2 port map( a => n3156, b => n3157, outb => n3155);
   U1933 : xor2 port map( a => n3159, b => n3160, outb => n3158);
   U1934 : xor2 port map( a => n3162, b => n3163, outb => n3161);
   U1935 : xor2 port map( a => n3165, b => n3166, outb => n3164);
   U1936 : xor2 port map( a => n3168, b => n3169, outb => n3167);
   U1937 : xor2 port map( a => n3170, b => n3171, outb => n282);
   U1938 : xor2 port map( a => mult_125_ab_1_12_port, b => 
                           mult_125_ab_0_13_port, outb => n3172);
   U1939 : xor2 port map( a => n3174, b => n3134, outb => n3173);
   U1940 : xor2 port map( a => n3176, b => n3177, outb => n3175);
   U1941 : xor2 port map( a => mult_125_ab_1_11_port, b => 
                           mult_125_ab_0_12_port, outb => n3178);
   U1942 : xor2 port map( a => n3180, b => n3172, outb => n3179);
   U1943 : xor2 port map( a => n3182, b => n3183, outb => n3181);
   U1944 : xor2 port map( a => n3185, b => n3186, outb => n3184);
   U1945 : xor2 port map( a => n3188, b => n3189, outb => n3187);
   U1946 : xor2 port map( a => n3191, b => n3192, outb => n3190);
   U1947 : xor2 port map( a => n3194, b => n3195, outb => n3193);
   U1948 : xor2 port map( a => n3197, b => n3198, outb => n3196);
   U1949 : xor2 port map( a => n3200, b => n3201, outb => n3199);
   U1950 : xor2 port map( a => n3203, b => n3204, outb => n3202);
   U1951 : xor2 port map( a => n3206, b => n3207, outb => n3205);
   U1952 : xor2 port map( a => n3209, b => n3210, outb => n3208);
   U1953 : xor2 port map( a => n3211, b => n3212, outb => n286);
   U1954 : xor2 port map( a => mult_125_ab_1_10_port, b => 
                           mult_125_ab_0_11_port, outb => n3213);
   U1955 : xor2 port map( a => n3215, b => n3178, outb => n3214);
   U1956 : xor2 port map( a => n3217, b => n3218, outb => n3216);
   U1957 : xor2 port map( a => n3220, b => n3221, outb => n3219);
   U1958 : xor2 port map( a => mult_125_ab_1_9_port, b => mult_125_ab_0_10_port
                           , outb => n3222);
   U1959 : xor2 port map( a => n3224, b => n3213, outb => n3223);
   U1960 : xor2 port map( a => n3226, b => n3227, outb => n3225);
   U1961 : xor2 port map( a => n3229, b => n3230, outb => n3228);
   U1962 : xor2 port map( a => n3232, b => n3233, outb => n3231);
   U1963 : xor2 port map( a => n3235, b => n3236, outb => n3234);
   U1964 : xor2 port map( a => n3238, b => n3239, outb => n3237);
   U1965 : xor2 port map( a => n3241, b => n3242, outb => n3240);
   U1966 : xor2 port map( a => n3244, b => n3245, outb => n3243);
   U1967 : xor2 port map( a => n3247, b => n3248, outb => n3246);
   U1968 : xor2 port map( a => n3250, b => n3251, outb => n3249);
   U1969 : xor2 port map( a => n3252, b => n3253, outb => n290);
   U1970 : xor2 port map( a => mult_125_ab_1_8_port, b => mult_125_ab_0_9_port,
                           outb => n3254);
   U1971 : xor2 port map( a => n3256, b => n3222, outb => n3255);
   U1972 : xor2 port map( a => n3258, b => n3259, outb => n3257);
   U1973 : xor2 port map( a => n3261, b => n3262, outb => n3260);
   U1974 : xor2 port map( a => n3264, b => n3265, outb => n3263);
   U1975 : xor2 port map( a => mult_125_ab_1_7_port, b => mult_125_ab_0_8_port,
                           outb => n3266);
   U1976 : xor2 port map( a => n3268, b => n3254, outb => n3267);
   U1977 : xor2 port map( a => n3270, b => n3271, outb => n3269);
   U1978 : xor2 port map( a => n3273, b => n3274, outb => n3272);
   U1979 : xor2 port map( a => n3276, b => n3277, outb => n3275);
   U1980 : xor2 port map( a => n3279, b => n3280, outb => n3278);
   U1981 : xor2 port map( a => n3282, b => n3283, outb => n3281);
   U1982 : xor2 port map( a => n3285, b => n3286, outb => n3284);
   U1983 : xor2 port map( a => n3288, b => n3289, outb => n3287);
   U1984 : xor2 port map( a => n3291, b => n3292, outb => n3290);
   U1985 : xor2 port map( a => n3293, b => n3294, outb => n294);
   U1986 : xor2 port map( a => mult_125_ab_1_6_port, b => mult_125_ab_0_7_port,
                           outb => n3295);
   U1987 : xor2 port map( a => n3297, b => n3266, outb => n3296);
   U1988 : xor2 port map( a => n3299, b => n3300, outb => n3298);
   U1989 : xor2 port map( a => n3302, b => n3303, outb => n3301);
   U1990 : xor2 port map( a => n3305, b => n3306, outb => n3304);
   U1991 : xor2 port map( a => n3308, b => n3309, outb => n3307);
   U1992 : xor2 port map( a => mult_125_ab_1_5_port, b => mult_125_ab_0_6_port,
                           outb => n3310);
   U1993 : xor2 port map( a => n3312, b => n3295, outb => n3311);
   U1994 : xor2 port map( a => n3314, b => n3315, outb => n3313);
   U1995 : xor2 port map( a => n3317, b => n3318, outb => n3316);
   U1996 : xor2 port map( a => n3320, b => n3321, outb => n3319);
   U1997 : xor2 port map( a => n3323, b => n3324, outb => n3322);
   U1998 : xor2 port map( a => n3326, b => n3327, outb => n3325);
   U1999 : xor2 port map( a => n3329, b => n3330, outb => n3328);
   U2000 : xor2 port map( a => n3332, b => n3333, outb => n3331);
   U2001 : xor2 port map( a => n3334, b => n3335, outb => n298);
   U2002 : xor2 port map( a => mult_125_ab_1_4_port, b => mult_125_ab_0_5_port,
                           outb => n3336);
   U2003 : xor2 port map( a => n3338, b => n3310, outb => n3337);
   U2004 : xor2 port map( a => n3340, b => n3341, outb => n3339);
   U2005 : xor2 port map( a => n3343, b => n3344, outb => n3342);
   U2006 : xor2 port map( a => n3346, b => n3347, outb => n3345);
   U2007 : xor2 port map( a => n3349, b => n3350, outb => n3348);
   U2008 : xor2 port map( a => n3352, b => n3353, outb => n3351);
   U2009 : xor2 port map( a => mult_125_ab_1_3_port, b => mult_125_ab_0_4_port,
                           outb => n3354);
   U2010 : xor2 port map( a => n3356, b => n3336, outb => n3355);
   U2011 : xor2 port map( a => n3358, b => n3359, outb => n3357);
   U2012 : xor2 port map( a => n3361, b => n3362, outb => n3360);
   U2013 : xor2 port map( a => n3364, b => n3365, outb => n3363);
   U2014 : xor2 port map( a => n3367, b => n3368, outb => n3366);
   U2015 : xor2 port map( a => n3370, b => n3371, outb => n3369);
   U2016 : xor2 port map( a => n3373, b => n3374, outb => n3372);
   U2017 : xor2 port map( a => n3375, b => n3376, outb => n303);
   U2018 : xor2 port map( a => mult_125_ab_1_2_port, b => mult_125_ab_0_3_port,
                           outb => n3377);
   U2019 : xor2 port map( a => n3379, b => n3354, outb => n3378);
   U2020 : xor2 port map( a => n3381, b => n3382, outb => n3380);
   U2021 : xor2 port map( a => n3384, b => n3385, outb => n3383);
   U2022 : xor2 port map( a => n3387, b => n3388, outb => n3386);
   U2023 : xor2 port map( a => n3390, b => n3391, outb => n3389);
   U2024 : xor2 port map( a => n3393, b => n3394, outb => n3392);
   U2025 : xor2 port map( a => n3396, b => n3397, outb => n3395);
   U2026 : xor2 port map( a => mult_125_ab_1_1_port, b => mult_125_ab_0_2_port,
                           outb => n3398);
   U2027 : xor2 port map( a => n3400, b => n3377, outb => n3399);
   U2028 : xor2 port map( a => n3402, b => n3403, outb => n3401);
   U2029 : xor2 port map( a => n3405, b => n3406, outb => n3404);
   U2030 : xor2 port map( a => n3408, b => n3409, outb => n3407);
   U2031 : xor2 port map( a => n3411, b => n3412, outb => n3410);
   U2032 : xor2 port map( a => n3414, b => n3415, outb => n3413);
   U2033 : xor2 port map( a => n3417, b => n3418, outb => n3416);
   U2034 : xor2 port map( a => n3419, b => n3410, outb => mult_125_A1_9_port);
   U2035 : xor2 port map( a => n3420, b => n3407, outb => mult_125_A1_7_port);
   U2036 : xor2 port map( a => n3421, b => n3404, outb => mult_125_A1_5_port);
   U2037 : xor2 port map( a => n3422, b => n3401, outb => mult_125_A1_3_port);
   U2038 : xor2 port map( a => n278, b => n277, outb => mult_125_A1_28_port);
   U2039 : xor2 port map( a => n282, b => n281, outb => mult_125_A1_26_port);
   U2040 : xor2 port map( a => n286, b => n285, outb => mult_125_A1_24_port);
   U2041 : xor2 port map( a => n290, b => n289, outb => mult_125_A1_22_port);
   U2042 : xor2 port map( a => n294, b => n293, outb => mult_125_A1_20_port);
   U2043 : xor2 port map( a => n3423, b => n3399, outb => mult_125_A1_1_port);
   U2044 : xor2 port map( a => n298, b => n297, outb => mult_125_A1_18_port);
   U2045 : xor2 port map( a => n303, b => n302, outb => mult_125_A1_16_port);
   U2046 : xor2 port map( a => n3424, b => n311, outb => mult_125_A1_13_port);
   U2047 : xor2 port map( a => n3425, b => n3413, outb => mult_125_A1_11_port);
   U2048 : xor2 port map( a => mult_125_G3_ab_1_0_port, b => 
                           mult_125_G3_ab_0_1_port, outb => n3426);
   U2049 : xor2 port map( a => n3427, b => n3428, outb => N99);
   U2050 : xor2 port map( a => n3429, b => n3430, outb => N98);
   U2051 : xor2 port map( a => n3431, b => n3432, outb => N97);
   U2052 : xor2 port map( a => n3433, b => n3434, outb => N96);
   U2053 : xor2 port map( a => n3435, b => n3436, outb => N95);
   U2054 : xor2 port map( a => n3437, b => n3438, outb => N94);
   U2055 : xor2 port map( a => n3439, b => n3440, outb => N93);
   U2056 : xor2 port map( a => n3441, b => n3442, outb => N92);
   U2057 : xor2 port map( a => n3443, b => n3444, outb => N91);
   U2058 : xor2 port map( a => n3445, b => n3446, outb => N90);
   U2059 : xor2 port map( a => mult_125_ab_1_0_port, b => mult_125_ab_0_1_port,
                           outb => n3447);
   U2060 : xor2 port map( a => n3448, b => n3449, outb => N9);
   U2061 : xor2 port map( a => n3450, b => n3451, outb => N89);
   U2062 : xor2 port map( a => n3452, b => n3453, outb => N88);
   U2063 : xor2 port map( a => n3454, b => n3455, outb => N87);
   U2064 : xor2 port map( a => n3456, b => n3457, outb => N86);
   U2065 : xor2 port map( a => n3458, b => n3459, outb => N85);
   U2066 : xor2 port map( a => n3460, b => n3461, outb => N84);
   U2067 : xor2 port map( a => n3462, b => n3463, outb => N83);
   U2068 : xor2 port map( a => n3464, b => n3465, outb => N82);
   U2069 : xor2 port map( a => n3466, b => n3467, outb => N81);
   U2070 : xor2 port map( a => n3468, b => n3469, outb => N80);
   U2071 : xor2 port map( a => n3470, b => n3471, outb => N8);
   U2072 : xor2 port map( a => n3472, b => n3473, outb => N79);
   U2073 : xor2 port map( a => n3474, b => n3475, outb => N78);
   U2074 : xor2 port map( a => n3476, b => n3477, outb => N77);
   U2075 : xor2 port map( a => n3478, b => n3479, outb => N76);
   U2076 : xor2 port map( a => n3480, b => n3481, outb => N75);
   U2077 : xor2 port map( a => n3482, b => n3483, outb => N74);
   U2078 : xor2 port map( a => mult_125_G2_ab_1_0_port, b => 
                           mult_125_G2_ab_0_1_port, outb => n3484);
   U2079 : xor2 port map( a => n3485, b => n2197, outb => N71);
   U2080 : xor2 port map( a => n2199, b => n3486, outb => N70);
   U2081 : xor2 port map( a => n3487, b => n3488, outb => N69);
   U2082 : xor2 port map( a => n3489, b => n3490, outb => N68);
   U2083 : xor2 port map( a => n3491, b => n3492, outb => N67);
   U2084 : xor2 port map( a => n3493, b => n3494, outb => N66);
   U2085 : xor2 port map( a => n3495, b => n3496, outb => N65);
   U2086 : xor2 port map( a => n3497, b => n3498, outb => N64);
   U2087 : xor2 port map( a => n3499, b => n3500, outb => N63);
   U2088 : xor2 port map( a => n3501, b => n3502, outb => N62);
   U2089 : xor2 port map( a => n3503, b => n3504, outb => N61);
   U2090 : xor2 port map( a => n3505, b => n3506, outb => N60);
   U2091 : xor2 port map( a => n3507, b => n3508, outb => N59);
   U2092 : xor2 port map( a => n3509, b => n3510, outb => N58);
   U2093 : xor2 port map( a => n3511, b => n3512, outb => N57);
   U2094 : xor2 port map( a => n3513, b => n3514, outb => N56);
   U2095 : xor2 port map( a => n3515, b => n3516, outb => N55);
   U2096 : xor2 port map( a => n3517, b => n3518, outb => N54);
   U2097 : xor2 port map( a => n3519, b => n3520, outb => N53);
   U2098 : xor2 port map( a => n3521, b => n3522, outb => N52);
   U2099 : xor2 port map( a => n3523, b => n3524, outb => N51);
   U2100 : xor2 port map( a => n3525, b => n3526, outb => N50);
   U2101 : xor2 port map( a => n3527, b => n3528, outb => N49);
   U2102 : xor2 port map( a => n3529, b => n3530, outb => N48);
   U2103 : xor2 port map( a => n3531, b => n3532, outb => N47);
   U2104 : xor2 port map( a => n3533, b => n3534, outb => N46);
   U2105 : xor2 port map( a => n3535, b => n3536, outb => N45);
   U2106 : xor2 port map( a => n3537, b => n3538, outb => N44);
   U2107 : xor2 port map( a => n3539, b => n3540, outb => N43);
   U2108 : xor2 port map( a => n3541, b => n3542, outb => N42);
   U2109 : xor2 port map( a => n3543, b => n3544, outb => N41);
   U2110 : xor2 port map( a => n3545, b => n2228, outb => N38);
   U2111 : xor2 port map( a => n2230, b => n3546, outb => N37);
   U2112 : xor2 port map( a => n3547, b => n3548, outb => N36);
   U2113 : xor2 port map( a => n3549, b => n3550, outb => N35);
   U2114 : xor2 port map( a => n3551, b => n3552, outb => N34);
   U2115 : xor2 port map( a => n3553, b => n3554, outb => N33);
   U2116 : xor2 port map( a => n3555, b => n3556, outb => N32);
   U2117 : xor2 port map( a => n3557, b => n3558, outb => N31);
   U2118 : xor2 port map( a => n3559, b => n3560, outb => N30);
   U2119 : xor2 port map( a => n3561, b => n3562, outb => N29);
   U2120 : xor2 port map( a => n3563, b => n3564, outb => N28);
   U2121 : xor2 port map( a => n3565, b => n3566, outb => N27);
   U2122 : xor2 port map( a => n3567, b => n3568, outb => N26);
   U2123 : xor2 port map( a => n3569, b => n3570, outb => N25);
   U2124 : xor2 port map( a => n3571, b => n3572, outb => N24);
   U2125 : xor2 port map( a => n3573, b => n3574, outb => N23);
   U2126 : xor2 port map( a => n3575, b => n3576, outb => N22);
   U2127 : xor2 port map( a => n3577, b => n3578, outb => N21);
   U2128 : xor2 port map( a => n3579, b => n3580, outb => N20);
   U2129 : xor2 port map( a => n3581, b => n3582, outb => N19);
   U2130 : xor2 port map( a => n3583, b => n3584, outb => N18);
   U2131 : xor2 port map( a => n3585, b => n3586, outb => N17);
   U2132 : xor2 port map( a => n3587, b => n3588, outb => N16);
   U2133 : xor2 port map( a => n3589, b => n3590, outb => N15);
   U2134 : xor2 port map( a => n3591, b => n3592, outb => N14);
   U2135 : xor2 port map( a => n3593, b => n3594, outb => N13);
   U2136 : xor2 port map( a => n3595, b => n3596, outb => N12);
   U2137 : xor2 port map( a => n3597, b => n3598, outb => N11);
   U2138 : xor2 port map( a => n3599, b => n2235, outb => N104);
   U2139 : xor2 port map( a => n2237, b => n3600, outb => N103);
   U2140 : xor2 port map( a => n3601, b => n3602, outb => N102);
   U2141 : xor2 port map( a => n3603, b => n3604, outb => N101);
   U2142 : xor2 port map( a => n3605, b => n3606, outb => N100);
   U2143 : xor2 port map( a => n3607, b => n3608, outb => N10);
   U2144 : nand2 port map( a => mult_125_G4_ab_0_15_port, b => 
                           mult_125_G4_ab_1_14_port, outb => n3609);
   U2145 : inv port map( inb => mult_125_G4_ab_3_15_port, outb => n3610);
   U2146 : inv port map( inb => mult_125_G4_ab_4_14_port, outb => n3611);
   U2147 : inv port map( inb => mult_125_G4_ab_5_15_port, outb => n3612);
   U2148 : inv port map( inb => mult_125_G4_ab_6_14_port, outb => n3613);
   U2149 : inv port map( inb => mult_125_G4_ab_7_15_port, outb => n3614);
   U2150 : inv port map( inb => mult_125_G4_ab_8_14_port, outb => n3615);
   U2151 : inv port map( inb => mult_125_G4_ab_9_15_port, outb => n3616);
   U2152 : inv port map( inb => mult_125_G4_ab_10_14_port, outb => n3617);
   U2153 : inv port map( inb => mult_125_G4_ab_11_15_port, outb => n3618);
   U2154 : inv port map( inb => mult_125_G4_ab_12_14_port, outb => n3619);
   U2155 : nand2 port map( a => mult_125_G4_ab_0_14_port, b => 
                           mult_125_G4_ab_1_13_port, outb => n400);
   U2156 : aoi22 port map( a => mult_125_G4_ab_2_13_port, b => n3620, c => n398
                           , d => n2240, outb => n403);
   U2157 : oai22 port map( a => n403, b => n402, c => n3621, d => n2241, outb 
                           => n405);
   U2158 : aoi22 port map( a => n405, b => mult_125_G4_ab_4_13_port, c => n3623
                           , d => n2248, outb => n3622);
   U2159 : oai22 port map( a => n3622, b => n3624, c => n406, d => n2251, outb 
                           => n409);
   U2160 : aoi22 port map( a => n409, b => mult_125_G4_ab_6_13_port, c => n3626
                           , d => n2254, outb => n3625);
   U2161 : inv port map( inb => mult_125_G4_ab_7_13_port, outb => n3627);
   U2162 : oai22 port map( a => n3625, b => n3627, c => n410, d => n2257, outb 
                           => n413);
   U2163 : aoi22 port map( a => n413, b => mult_125_G4_ab_8_13_port, c => n3629
                           , d => n2260, outb => n3628);
   U2164 : inv port map( inb => mult_125_G4_ab_9_13_port, outb => n3630);
   U2165 : oai22 port map( a => n3628, b => n3630, c => n414, d => n2263, outb 
                           => n417);
   U2166 : aoi22 port map( a => n417, b => mult_125_G4_ab_10_13_port, c => 
                           n3632, d => n2266, outb => n3631);
   U2167 : inv port map( inb => mult_125_G4_ab_11_13_port, outb => n3633);
   U2168 : oai22 port map( a => n3631, b => n3633, c => n418, d => n2269, outb 
                           => n421);
   U2169 : aoi22 port map( a => n421, b => mult_125_G4_ab_12_13_port, c => 
                           n3635, d => n2272, outb => n3634);
   U2170 : inv port map( inb => mult_125_G4_ab_13_13_port, outb => n3636);
   U2171 : oai22 port map( a => n3634, b => n3636, c => n422, d => n2275, outb 
                           => n425);
   U2172 : aoi22 port map( a => n425, b => mult_125_G4_ab_14_13_port, c => 
                           n3638, d => n2278, outb => n3637);
   U2173 : nand2 port map( a => mult_125_G4_ab_0_13_port, b => 
                           mult_125_G4_ab_1_12_port, outb => n430);
   U2174 : aoi22 port map( a => mult_125_G4_ab_2_12_port, b => n3640, c => n428
                           , d => n2243, outb => n3639);
   U2175 : oai22 port map( a => n3639, b => n3641, c => n431, d => n2244, outb 
                           => n434);
   U2176 : aoi22 port map( a => n434, b => mult_125_G4_ab_4_12_port, c => n3643
                           , d => n2286, outb => n3642);
   U2177 : aoi22 port map( a => n436, b => mult_125_G4_ab_5_12_port, c => n3645
                           , d => n2246, outb => n3644);
   U2178 : inv port map( inb => mult_125_G4_ab_6_12_port, outb => n3646);
   U2179 : oai22 port map( a => n3644, b => n3646, c => n437, d => n2249, outb 
                           => n440);
   U2180 : aoi22 port map( a => n440, b => mult_125_G4_ab_7_12_port, c => n3648
                           , d => n2252, outb => n3647);
   U2181 : inv port map( inb => mult_125_G4_ab_8_12_port, outb => n3649);
   U2182 : oai22 port map( a => n3647, b => n3649, c => n441, d => n2255, outb 
                           => n444);
   U2183 : aoi22 port map( a => n444, b => mult_125_G4_ab_9_12_port, c => n3651
                           , d => n2258, outb => n3650);
   U2184 : inv port map( inb => mult_125_G4_ab_10_12_port, outb => n3652);
   U2185 : oai22 port map( a => n3650, b => n3652, c => n445, d => n2261, outb 
                           => n448);
   U2186 : aoi22 port map( a => n448, b => mult_125_G4_ab_11_12_port, c => 
                           n3654, d => n2264, outb => n3653);
   U2187 : inv port map( inb => mult_125_G4_ab_12_12_port, outb => n3655);
   U2188 : oai22 port map( a => n3653, b => n3655, c => n449, d => n2267, outb 
                           => n452);
   U2189 : aoi22 port map( a => n452, b => mult_125_G4_ab_13_12_port, c => 
                           n3657, d => n2270, outb => n3656);
   U2190 : inv port map( inb => mult_125_G4_ab_14_12_port, outb => n3658);
   U2191 : oai22 port map( a => n3656, b => n3658, c => n453, d => n2273, outb 
                           => n456);
   U2192 : nand2 port map( a => mult_125_G4_ab_0_12_port, b => 
                           mult_125_G4_ab_1_11_port, outb => n459);
   U2193 : aoi22 port map( a => mult_125_G4_ab_2_11_port, b => n3659, c => n457
                           , d => n2281, outb => n462);
   U2194 : oai22 port map( a => n462, b => n461, c => n3660, d => n2282, outb 
                           => n464);
   U2195 : oai22 port map( a => n3661, b => n3662, c => n463, d => n2292, outb 
                           => n466);
   U2196 : aoi22 port map( a => n466, b => mult_125_G4_ab_5_11_port, c => n3664
                           , d => n2284, outb => n3663);
   U2197 : oai22 port map( a => n3663, b => n3665, c => n467, d => n2295, outb 
                           => n470);
   U2198 : oai22 port map( a => n3666, b => n3667, c => n469, d => n2298, outb 
                           => n472);
   U2199 : aoi22 port map( a => n472, b => mult_125_G4_ab_8_11_port, c => n3669
                           , d => n2301, outb => n3668);
   U2200 : inv port map( inb => mult_125_G4_ab_9_11_port, outb => n3670);
   U2201 : oai22 port map( a => n3668, b => n3670, c => n473, d => n2304, outb 
                           => n476);
   U2202 : aoi22 port map( a => n476, b => mult_125_G4_ab_10_11_port, c => 
                           n3672, d => n2307, outb => n3671);
   U2203 : inv port map( inb => mult_125_G4_ab_11_11_port, outb => n3673);
   U2204 : oai22 port map( a => n3671, b => n3673, c => n477, d => n2310, outb 
                           => n480);
   U2205 : aoi22 port map( a => n480, b => mult_125_G4_ab_12_11_port, c => 
                           n3675, d => n2313, outb => n3674);
   U2206 : inv port map( inb => mult_125_G4_ab_13_11_port, outb => n3676);
   U2207 : oai22 port map( a => n3674, b => n3676, c => n481, d => n2316, outb 
                           => n484);
   U2208 : aoi22 port map( a => n484, b => mult_125_G4_ab_14_11_port, c => 
                           n3677, d => n2319, outb => n487);
   U2209 : nand2 port map( a => mult_125_G4_ab_0_11_port, b => 
                           mult_125_G4_ab_1_10_port, outb => n490);
   U2210 : aoi22 port map( a => mult_125_G4_ab_2_10_port, b => n3679, c => n488
                           , d => n2287, outb => n3678);
   U2211 : oai22 port map( a => n3678, b => n3680, c => n491, d => n2288, outb 
                           => n494);
   U2212 : aoi22 port map( a => n494, b => mult_125_G4_ab_4_10_port, c => n3681
                           , d => n2327, outb => n497);
   U2213 : oai22 port map( a => n497, b => n496, c => n3682, d => n2290, outb 
                           => n499);
   U2214 : aoi22 port map( a => n499, b => mult_125_G4_ab_6_10_port, c => n3684
                           , d => n2330, outb => n3683);
   U2215 : oai22 port map( a => n3683, b => n3685, c => n500, d => n2293, outb 
                           => n503);
   U2216 : inv port map( inb => mult_125_G4_ab_8_10_port, outb => n3686);
   U2217 : oai22 port map( a => n3687, b => n3686, c => n502, d => n2296, outb 
                           => n505);
   U2218 : aoi22 port map( a => n505, b => mult_125_G4_ab_9_10_port, c => n3689
                           , d => n2299, outb => n3688);
   U2219 : inv port map( inb => mult_125_G4_ab_10_10_port, outb => n3690);
   U2220 : oai22 port map( a => n3688, b => n3690, c => n506, d => n2302, outb 
                           => n509);
   U2221 : aoi22 port map( a => n509, b => mult_125_G4_ab_11_10_port, c => 
                           n3692, d => n2305, outb => n3691);
   U2222 : inv port map( inb => mult_125_G4_ab_12_10_port, outb => n3693);
   U2223 : oai22 port map( a => n3691, b => n3693, c => n510, d => n2308, outb 
                           => n513);
   U2224 : aoi22 port map( a => n513, b => mult_125_G4_ab_13_10_port, c => 
                           n3695, d => n2311, outb => n3694);
   U2225 : inv port map( inb => mult_125_G4_ab_14_10_port, outb => n3696);
   U2226 : oai22 port map( a => n3694, b => n3696, c => n514, d => n2314, outb 
                           => n517);
   U2227 : nand2 port map( a => mult_125_G4_ab_0_10_port, b => 
                           mult_125_G4_ab_1_9_port, outb => n520);
   U2228 : aoi22 port map( a => mult_125_G4_ab_2_9_port, b => n3698, c => n518,
                           d => n2322, outb => n3697);
   U2229 : oai22 port map( a => n3697, b => n3699, c => n521, d => n2323, outb 
                           => n524);
   U2230 : oai22 port map( a => n3700, b => n3701, c => n523, d => n2336, outb 
                           => n526);
   U2231 : aoi22 port map( a => n526, b => mult_125_G4_ab_5_9_port, c => n3703,
                           d => n2325, outb => n3702);
   U2232 : oai22 port map( a => n3702, b => n3704, c => n527, d => n2339, outb 
                           => n530);
   U2233 : aoi22 port map( a => n530, b => mult_125_G4_ab_7_9_port, c => n3706,
                           d => n2328, outb => n3705);
   U2234 : oai22 port map( a => n3705, b => n3707, c => n531, d => n2342, outb 
                           => n534);
   U2235 : oai22 port map( a => n3708, b => n3709, c => n533, d => n2345, outb 
                           => n536);
   U2236 : aoi22 port map( a => n536, b => mult_125_G4_ab_10_9_port, c => n3711
                           , d => n2348, outb => n3710);
   U2237 : inv port map( inb => mult_125_G4_ab_11_9_port, outb => n3712);
   U2238 : oai22 port map( a => n3710, b => n3712, c => n537, d => n2351, outb 
                           => n540);
   U2239 : aoi22 port map( a => n540, b => mult_125_G4_ab_12_9_port, c => n3714
                           , d => n2354, outb => n3713);
   U2240 : inv port map( inb => mult_125_G4_ab_13_9_port, outb => n3715);
   U2241 : oai22 port map( a => n3713, b => n3715, c => n541, d => n2357, outb 
                           => n544);
   U2242 : aoi22 port map( a => n544, b => mult_125_G4_ab_14_9_port, c => n3716
                           , d => n2360, outb => n547);
   U2243 : nand2 port map( a => mult_125_G4_ab_0_9_port, b => 
                           mult_125_G4_ab_1_8_port, outb => n550);
   U2244 : aoi22 port map( a => mult_125_G4_ab_2_8_port, b => n3718, c => n548,
                           d => n2331, outb => n3717);
   U2245 : oai22 port map( a => n3717, b => n3719, c => n551, d => n2332, outb 
                           => n554);
   U2246 : oai22 port map( a => n3720, b => n3721, c => n553, d => n2368, outb 
                           => n556);
   U2247 : oai22 port map( a => n3722, b => n3723, c => n555, d => n2334, outb 
                           => n558);
   U2248 : aoi22 port map( a => n558, b => mult_125_G4_ab_6_8_port, c => n3725,
                           d => n2371, outb => n3724);
   U2249 : oai22 port map( a => n3724, b => n3726, c => n559, d => n2337, outb 
                           => n562);
   U2250 : aoi22 port map( a => n562, b => mult_125_G4_ab_8_8_port, c => n3728,
                           d => n2374, outb => n3727);
   U2251 : oai22 port map( a => n3727, b => n3729, c => n563, d => n2340, outb 
                           => n566);
   U2252 : inv port map( inb => mult_125_G4_ab_10_8_port, outb => n3730);
   U2253 : oai22 port map( a => n3731, b => n3730, c => n565, d => n2343, outb 
                           => n568);
   U2254 : aoi22 port map( a => n568, b => mult_125_G4_ab_11_8_port, c => n3733
                           , d => n2346, outb => n3732);
   U2255 : inv port map( inb => mult_125_G4_ab_12_8_port, outb => n3734);
   U2256 : oai22 port map( a => n3732, b => n3734, c => n569, d => n2349, outb 
                           => n572);
   U2257 : aoi22 port map( a => n572, b => mult_125_G4_ab_13_8_port, c => n3736
                           , d => n2352, outb => n3735);
   U2258 : inv port map( inb => mult_125_G4_ab_14_8_port, outb => n3737);
   U2259 : oai22 port map( a => n3735, b => n3737, c => n573, d => n2355, outb 
                           => n576);
   U2260 : nand2 port map( a => mult_125_G4_ab_0_8_port, b => 
                           mult_125_G4_ab_1_7_port, outb => n579);
   U2261 : aoi22 port map( a => mult_125_G4_ab_2_7_port, b => n3738, c => n577,
                           d => n2363, outb => n582);
   U2262 : oai22 port map( a => n582, b => n581, c => n3739, d => n2364, outb 
                           => n584);
   U2263 : oai22 port map( a => n3740, b => n3741, c => n583, d => n2380, outb 
                           => n586);
   U2264 : aoi22 port map( a => n586, b => mult_125_G4_ab_5_7_port, c => n3743,
                           d => n2366, outb => n3742);
   U2265 : oai22 port map( a => n3742, b => n3744, c => n587, d => n2383, outb 
                           => n590);
   U2266 : aoi22 port map( a => n590, b => mult_125_G4_ab_7_7_port, c => n3746,
                           d => n2369, outb => n3745);
   U2267 : oai22 port map( a => n3745, b => n3747, c => n591, d => n2386, outb 
                           => n594);
   U2268 : aoi22 port map( a => n594, b => mult_125_G4_ab_9_7_port, c => n3749,
                           d => n2372, outb => n3748);
   U2269 : oai22 port map( a => n3748, b => n3750, c => n595, d => n2389, outb 
                           => n598);
   U2270 : oai22 port map( a => n3751, b => n3752, c => n597, d => n2392, outb 
                           => n600);
   U2271 : aoi22 port map( a => n600, b => mult_125_G4_ab_12_7_port, c => n3754
                           , d => n2395, outb => n3753);
   U2272 : inv port map( inb => mult_125_G4_ab_13_7_port, outb => n3755);
   U2273 : oai22 port map( a => n3753, b => n3755, c => n601, d => n2398, outb 
                           => n604);
   U2274 : aoi22 port map( a => n604, b => mult_125_G4_ab_14_7_port, c => n3756
                           , d => n2401, outb => n607);
   U2275 : nand2 port map( a => mult_125_G4_ab_0_7_port, b => 
                           mult_125_G4_ab_1_6_port, outb => n610);
   U2276 : aoi22 port map( a => mult_125_G4_ab_2_6_port, b => n3758, c => n608,
                           d => n2375, outb => n3757);
   U2277 : oai22 port map( a => n3757, b => n3759, c => n611, d => n2376, outb 
                           => n614);
   U2278 : aoi22 port map( a => n614, b => mult_125_G4_ab_4_6_port, c => n3760,
                           d => n2409, outb => n617);
   U2279 : oai22 port map( a => n617, b => n616, c => n3761, d => n2378, outb 
                           => n619);
   U2280 : aoi22 port map( a => n619, b => mult_125_G4_ab_6_6_port, c => n3763,
                           d => n2412, outb => n3762);
   U2281 : oai22 port map( a => n3762, b => n3764, c => n620, d => n2381, outb 
                           => n623);
   U2282 : aoi22 port map( a => n623, b => mult_125_G4_ab_8_6_port, c => n3765,
                           d => n2415, outb => n626);
   U2283 : oai22 port map( a => n626, b => n625, c => n3766, d => n2384, outb 
                           => n628);
   U2284 : aoi22 port map( a => n628, b => mult_125_G4_ab_10_6_port, c => n3768
                           , d => n2418, outb => n3767);
   U2285 : oai22 port map( a => n3767, b => n3769, c => n629, d => n2387, outb 
                           => n632);
   U2286 : inv port map( inb => mult_125_G4_ab_12_6_port, outb => n3770);
   U2287 : oai22 port map( a => n3771, b => n3770, c => n631, d => n2390, outb 
                           => n634);
   U2288 : aoi22 port map( a => n634, b => mult_125_G4_ab_13_6_port, c => n3773
                           , d => n2393, outb => n3772);
   U2289 : inv port map( inb => mult_125_G4_ab_14_6_port, outb => n3774);
   U2290 : oai22 port map( a => n3772, b => n3774, c => n635, d => n2396, outb 
                           => n638);
   U2291 : nand2 port map( a => mult_125_G4_ab_0_6_port, b => 
                           mult_125_G4_ab_1_5_port, outb => n641);
   U2292 : aoi22 port map( a => mult_125_G4_ab_2_5_port, b => n3775, c => n639,
                           d => n2404, outb => n644);
   U2293 : oai22 port map( a => n644, b => n643, c => n3776, d => n2405, outb 
                           => n646);
   U2294 : oai22 port map( a => n3777, b => n3778, c => n645, d => n2424, outb 
                           => n648);
   U2295 : aoi22 port map( a => n648, b => mult_125_G4_ab_5_5_port, c => n3779,
                           d => n2407, outb => n651);
   U2296 : oai22 port map( a => n651, b => n650, c => n3780, d => n2427, outb 
                           => n653);
   U2297 : aoi22 port map( a => n653, b => mult_125_G4_ab_7_5_port, c => n3782,
                           d => n2410, outb => n3781);
   U2298 : oai22 port map( a => n3781, b => n3783, c => n654, d => n2430, outb 
                           => n657);
   U2299 : aoi22 port map( a => n657, b => mult_125_G4_ab_9_5_port, c => n3785,
                           d => n2413, outb => n3784);
   U2300 : oai22 port map( a => n3784, b => n3786, c => n658, d => n2433, outb 
                           => n661);
   U2301 : aoi22 port map( a => n661, b => mult_125_G4_ab_11_5_port, c => n3788
                           , d => n2416, outb => n3787);
   U2302 : oai22 port map( a => n3787, b => n3789, c => n662, d => n2436, outb 
                           => n665);
   U2303 : oai22 port map( a => n3790, b => n3791, c => n664, d => n2439, outb 
                           => n667);
   U2304 : aoi22 port map( a => n667, b => mult_125_G4_ab_14_5_port, c => n3792
                           , d => n2442, outb => n670);
   U2305 : nand2 port map( a => mult_125_G4_ab_0_5_port, b => 
                           mult_125_G4_ab_1_4_port, outb => n673);
   U2306 : aoi22 port map( a => mult_125_G4_ab_2_4_port, b => n3794, c => n671,
                           d => n2419, outb => n3793);
   U2307 : oai22 port map( a => n3793, b => n3795, c => n674, d => n2420, outb 
                           => n677);
   U2308 : aoi22 port map( a => n677, b => mult_125_G4_ab_4_4_port, c => n3796,
                           d => n2450, outb => n680);
   U2309 : oai22 port map( a => n680, b => n679, c => n3797, d => n2422, outb 
                           => n682);
   U2310 : aoi22 port map( a => n682, b => mult_125_G4_ab_6_4_port, c => n3798,
                           d => n2453, outb => n685);
   U2311 : oai22 port map( a => n685, b => n684, c => n3799, d => n2425, outb 
                           => n687);
   U2312 : aoi22 port map( a => n687, b => mult_125_G4_ab_8_4_port, c => n3801,
                           d => n2456, outb => n3800);
   U2313 : oai22 port map( a => n3800, b => n3802, c => n688, d => n2428, outb 
                           => n691);
   U2314 : aoi22 port map( a => n691, b => mult_125_G4_ab_10_4_port, c => n3803
                           , d => n2459, outb => n694);
   U2315 : oai22 port map( a => n694, b => n693, c => n3804, d => n2431, outb 
                           => n696);
   U2316 : aoi22 port map( a => n696, b => mult_125_G4_ab_12_4_port, c => n3806
                           , d => n2462, outb => n3805);
   U2317 : oai22 port map( a => n3805, b => n3807, c => n697, d => n2434, outb 
                           => n700);
   U2318 : aoi22 port map( a => n700, b => mult_125_G4_ab_14_4_port, c => n3808
                           , d => n2437, outb => n703);
   U2319 : nand2 port map( a => mult_125_G4_ab_0_4_port, b => 
                           mult_125_G4_ab_1_3_port, outb => n706);
   U2320 : aoi22 port map( a => mult_125_G4_ab_2_3_port, b => n3809, c => n704,
                           d => n2445, outb => n709);
   U2321 : oai22 port map( a => n709, b => n708, c => n3810, d => n2446, outb 
                           => n711);
   U2322 : oai22 port map( a => n3811, b => n3812, c => n710, d => n2468, outb 
                           => n713);
   U2323 : aoi22 port map( a => n713, b => mult_125_G4_ab_5_3_port, c => n3814,
                           d => n2448, outb => n3813);
   U2324 : oai22 port map( a => n3813, b => n3815, c => n714, d => n2471, outb 
                           => n717);
   U2325 : aoi22 port map( a => n717, b => mult_125_G4_ab_7_3_port, c => n3817,
                           d => n2451, outb => n3816);
   U2326 : oai22 port map( a => n3816, b => n3818, c => n718, d => n2474, outb 
                           => n721);
   U2327 : aoi22 port map( a => n721, b => mult_125_G4_ab_9_3_port, c => n3820,
                           d => n2454, outb => n3819);
   U2328 : oai22 port map( a => n3819, b => n3821, c => n722, d => n2477, outb 
                           => n725);
   U2329 : aoi22 port map( a => n725, b => mult_125_G4_ab_11_3_port, c => n3823
                           , d => n2457, outb => n3822);
   U2330 : oai22 port map( a => n3822, b => n3824, c => n726, d => n2480, outb 
                           => n729);
   U2331 : aoi22 port map( a => n729, b => mult_125_G4_ab_13_3_port, c => n3826
                           , d => n2460, outb => n3825);
   U2332 : inv port map( inb => mult_125_G4_ab_14_3_port, outb => n3827);
   U2333 : oai22 port map( a => n3825, b => n3827, c => n730, d => n2483, outb 
                           => n733);
   U2334 : nand2 port map( a => mult_125_G4_ab_0_3_port, b => 
                           mult_125_G4_ab_1_2_port, outb => n736);
   U2335 : aoi22 port map( a => mult_125_G4_ab_2_2_port, b => n3829, c => n734,
                           d => n2463, outb => n3828);
   U2336 : oai22 port map( a => n3828, b => n3830, c => n737, d => n2464, outb 
                           => n740);
   U2337 : aoi22 port map( a => n740, b => mult_125_G4_ab_4_2_port, c => n3832,
                           d => n2491, outb => n3831);
   U2338 : oai22 port map( a => n3831, b => n3833, c => n741, d => n2466, outb 
                           => n744);
   U2339 : aoi22 port map( a => n744, b => mult_125_G4_ab_6_2_port, c => n3834,
                           d => n2494, outb => n747);
   U2340 : oai22 port map( a => n747, b => n746, c => n3835, d => n2469, outb 
                           => n749);
   U2341 : aoi22 port map( a => n749, b => mult_125_G4_ab_8_2_port, c => n3837,
                           d => n2497, outb => n3836);
   U2342 : oai22 port map( a => n3836, b => n3838, c => n750, d => n2472, outb 
                           => n753);
   U2343 : aoi22 port map( a => n753, b => mult_125_G4_ab_10_2_port, c => n3840
                           , d => n2500, outb => n3839);
   U2344 : oai22 port map( a => n3839, b => n3841, c => n754, d => n2475, outb 
                           => n757);
   U2345 : aoi22 port map( a => n757, b => mult_125_G4_ab_12_2_port, c => n3843
                           , d => n2503, outb => n3842);
   U2346 : oai22 port map( a => n3842, b => n3844, c => n758, d => n2478, outb 
                           => n761);
   U2347 : aoi22 port map( a => n761, b => mult_125_G4_ab_14_2_port, c => n3846
                           , d => n2506, outb => n3845);
   U2348 : nand2 port map( a => mult_125_G4_ab_0_2_port, b => 
                           mult_125_G4_ab_1_1_port, outb => n766);
   U2349 : aoi22 port map( a => mult_125_G4_ab_2_1_port, b => n3848, c => n764,
                           d => n2486, outb => n3847);
   U2350 : oai22 port map( a => n3847, b => n3849, c => n767, d => n2487, outb 
                           => n770);
   U2351 : inv port map( inb => mult_125_G4_ab_4_1_port, outb => n3850);
   U2352 : oai22 port map( a => n3851, b => n3850, c => n769, d => n2512, outb 
                           => n772);
   U2353 : aoi22 port map( a => n772, b => mult_125_G4_ab_5_1_port, c => n3853,
                           d => n2489, outb => n3852);
   U2354 : oai22 port map( a => n3852, b => n3854, c => n773, d => n2515, outb 
                           => n776);
   U2355 : aoi22 port map( a => n776, b => mult_125_G4_ab_7_1_port, c => n3856,
                           d => n2492, outb => n3855);
   U2356 : oai22 port map( a => n3855, b => n3857, c => n777, d => n2518, outb 
                           => n780);
   U2357 : aoi22 port map( a => n780, b => mult_125_G4_ab_9_1_port, c => n3859,
                           d => n2495, outb => n3858);
   U2358 : oai22 port map( a => n3858, b => n3860, c => n781, d => n2521, outb 
                           => n784);
   U2359 : aoi22 port map( a => n784, b => mult_125_G4_ab_11_1_port, c => n3862
                           , d => n2498, outb => n3861);
   U2360 : oai22 port map( a => n3861, b => n3863, c => n785, d => n2524, outb 
                           => n788);
   U2361 : aoi22 port map( a => n788, b => mult_125_G4_ab_13_1_port, c => n3865
                           , d => n2501, outb => n3864);
   U2362 : inv port map( inb => mult_125_G4_ab_14_1_port, outb => n3866);
   U2363 : oai22 port map( a => n3864, b => n3866, c => n789, d => n2527, outb 
                           => n792);
   U2364 : nand2 port map( a => mult_125_G4_ab_1_0_port, b => 
                           mult_125_G4_ab_0_1_port, outb => n3867);
   U2365 : aoi22 port map( a => mult_125_G4_ab_2_0_port, b => n794, c => n3869,
                           d => n2507, outb => n3868);
   U2366 : aoi22 port map( a => n796, b => mult_125_G4_ab_3_0_port, c => n3871,
                           d => n2508, outb => n3870);
   U2367 : inv port map( inb => mult_125_G4_ab_4_0_port, outb => n3872);
   U2368 : oai22 port map( a => n3870, b => n3872, c => n797, d => n3873, outb 
                           => n800);
   U2369 : aoi22 port map( a => n800, b => mult_125_G4_ab_5_0_port, c => n3875,
                           d => n2510, outb => n3874);
   U2370 : inv port map( inb => mult_125_G4_ab_6_0_port, outb => n3876);
   U2371 : oai22 port map( a => n3874, b => n3876, c => n801, d => n3877, outb 
                           => n804);
   U2372 : aoi22 port map( a => n804, b => mult_125_G4_ab_7_0_port, c => n3879,
                           d => n2513, outb => n3878);
   U2373 : inv port map( inb => mult_125_G4_ab_8_0_port, outb => n3880);
   U2374 : oai22 port map( a => n3878, b => n3880, c => n805, d => n3881, outb 
                           => n808);
   U2375 : aoi22 port map( a => n808, b => mult_125_G4_ab_9_0_port, c => n3883,
                           d => n2516, outb => n3882);
   U2376 : inv port map( inb => mult_125_G4_ab_10_0_port, outb => n3884);
   U2377 : oai22 port map( a => n3882, b => n3884, c => n809, d => n3885, outb 
                           => n812);
   U2378 : aoi22 port map( a => n812, b => mult_125_G4_ab_11_0_port, c => n3887
                           , d => n2519, outb => n3886);
   U2379 : inv port map( inb => mult_125_G4_ab_12_0_port, outb => n3888);
   U2380 : oai22 port map( a => n3886, b => n3888, c => n813, d => n3889, outb 
                           => n816);
   U2381 : aoi22 port map( a => n816, b => mult_125_G4_ab_13_0_port, c => n3891
                           , d => n2522, outb => n3890);
   U2382 : inv port map( inb => mult_125_G4_ab_14_0_port, outb => n3892);
   U2383 : oai22 port map( a => n3890, b => n3892, c => n817, d => n3893, outb 
                           => n820);
   U2384 : inv port map( inb => mult_125_G4_ZB, outb => n272);
   U2385 : inv port map( inb => mult_125_G4_ZA, outb => n273);
   U2386 : nand2 port map( a => mult_125_G3_ab_0_15_port, b => 
                           mult_125_G3_ab_1_14_port, outb => n3894);
   U2387 : inv port map( inb => mult_125_G3_ab_3_15_port, outb => n3895);
   U2388 : inv port map( inb => mult_125_G3_ab_4_14_port, outb => n3896);
   U2389 : inv port map( inb => mult_125_G3_ab_5_15_port, outb => n3897);
   U2390 : inv port map( inb => mult_125_G3_ab_6_14_port, outb => n3898);
   U2391 : inv port map( inb => mult_125_G3_ab_7_15_port, outb => n3899);
   U2392 : inv port map( inb => mult_125_G3_ab_8_14_port, outb => n3900);
   U2393 : inv port map( inb => mult_125_G3_ab_9_15_port, outb => n3901);
   U2394 : inv port map( inb => mult_125_G3_ab_10_14_port, outb => n3902);
   U2395 : inv port map( inb => mult_125_G3_ab_11_15_port, outb => n3903);
   U2396 : inv port map( inb => mult_125_G3_ab_12_14_port, outb => n3904);
   U2397 : nand2 port map( a => mult_125_G3_ab_0_14_port, b => 
                           mult_125_G3_ab_1_13_port, outb => n838);
   U2398 : aoi22 port map( a => mult_125_G3_ab_2_13_port, b => n3905, c => n836
                           , d => n2537, outb => n841);
   U2399 : oai22 port map( a => n841, b => n840, c => n3906, d => n2538, outb 
                           => n843);
   U2400 : aoi22 port map( a => n843, b => mult_125_G3_ab_4_13_port, c => n3908
                           , d => n2545, outb => n3907);
   U2401 : oai22 port map( a => n3907, b => n3909, c => n844, d => n2548, outb 
                           => n847);
   U2402 : aoi22 port map( a => n847, b => mult_125_G3_ab_6_13_port, c => n3911
                           , d => n2551, outb => n3910);
   U2403 : inv port map( inb => mult_125_G3_ab_7_13_port, outb => n3912);
   U2404 : oai22 port map( a => n3910, b => n3912, c => n848, d => n2554, outb 
                           => n851);
   U2405 : aoi22 port map( a => n851, b => mult_125_G3_ab_8_13_port, c => n3914
                           , d => n2557, outb => n3913);
   U2406 : inv port map( inb => mult_125_G3_ab_9_13_port, outb => n3915);
   U2407 : oai22 port map( a => n3913, b => n3915, c => n852, d => n2560, outb 
                           => n855);
   U2408 : aoi22 port map( a => n855, b => mult_125_G3_ab_10_13_port, c => 
                           n3917, d => n2563, outb => n3916);
   U2409 : inv port map( inb => mult_125_G3_ab_11_13_port, outb => n3918);
   U2410 : oai22 port map( a => n3916, b => n3918, c => n856, d => n2566, outb 
                           => n859);
   U2411 : aoi22 port map( a => n859, b => mult_125_G3_ab_12_13_port, c => 
                           n3920, d => n2569, outb => n3919);
   U2412 : inv port map( inb => mult_125_G3_ab_13_13_port, outb => n3921);
   U2413 : oai22 port map( a => n3919, b => n3921, c => n860, d => n2572, outb 
                           => n863);
   U2414 : aoi22 port map( a => n863, b => mult_125_G3_ab_14_13_port, c => 
                           n3923, d => n2575, outb => n3922);
   U2415 : nand2 port map( a => mult_125_G3_ab_0_13_port, b => 
                           mult_125_G3_ab_1_12_port, outb => n868);
   U2416 : aoi22 port map( a => mult_125_G3_ab_2_12_port, b => n3925, c => n866
                           , d => n2540, outb => n3924);
   U2417 : oai22 port map( a => n3924, b => n3926, c => n869, d => n2541, outb 
                           => n872);
   U2418 : aoi22 port map( a => n872, b => mult_125_G3_ab_4_12_port, c => n3928
                           , d => n2583, outb => n3927);
   U2419 : aoi22 port map( a => n874, b => mult_125_G3_ab_5_12_port, c => n3930
                           , d => n2543, outb => n3929);
   U2420 : inv port map( inb => mult_125_G3_ab_6_12_port, outb => n3931);
   U2421 : oai22 port map( a => n3929, b => n3931, c => n875, d => n2546, outb 
                           => n878);
   U2422 : aoi22 port map( a => n878, b => mult_125_G3_ab_7_12_port, c => n3933
                           , d => n2549, outb => n3932);
   U2423 : inv port map( inb => mult_125_G3_ab_8_12_port, outb => n3934);
   U2424 : oai22 port map( a => n3932, b => n3934, c => n879, d => n2552, outb 
                           => n882);
   U2425 : aoi22 port map( a => n882, b => mult_125_G3_ab_9_12_port, c => n3936
                           , d => n2555, outb => n3935);
   U2426 : inv port map( inb => mult_125_G3_ab_10_12_port, outb => n3937);
   U2427 : oai22 port map( a => n3935, b => n3937, c => n883, d => n2558, outb 
                           => n886);
   U2428 : aoi22 port map( a => n886, b => mult_125_G3_ab_11_12_port, c => 
                           n3939, d => n2561, outb => n3938);
   U2429 : inv port map( inb => mult_125_G3_ab_12_12_port, outb => n3940);
   U2430 : oai22 port map( a => n3938, b => n3940, c => n887, d => n2564, outb 
                           => n890);
   U2431 : aoi22 port map( a => n890, b => mult_125_G3_ab_13_12_port, c => 
                           n3942, d => n2567, outb => n3941);
   U2432 : inv port map( inb => mult_125_G3_ab_14_12_port, outb => n3943);
   U2433 : oai22 port map( a => n3941, b => n3943, c => n891, d => n2570, outb 
                           => n894);
   U2434 : nand2 port map( a => mult_125_G3_ab_0_12_port, b => 
                           mult_125_G3_ab_1_11_port, outb => n897);
   U2435 : aoi22 port map( a => mult_125_G3_ab_2_11_port, b => n3944, c => n895
                           , d => n2578, outb => n900);
   U2436 : oai22 port map( a => n900, b => n899, c => n3945, d => n2579, outb 
                           => n902);
   U2437 : oai22 port map( a => n3946, b => n3947, c => n901, d => n2589, outb 
                           => n904);
   U2438 : aoi22 port map( a => n904, b => mult_125_G3_ab_5_11_port, c => n3949
                           , d => n2581, outb => n3948);
   U2439 : oai22 port map( a => n3948, b => n3950, c => n905, d => n2592, outb 
                           => n908);
   U2440 : oai22 port map( a => n3951, b => n3952, c => n907, d => n2595, outb 
                           => n910);
   U2441 : aoi22 port map( a => n910, b => mult_125_G3_ab_8_11_port, c => n3954
                           , d => n2598, outb => n3953);
   U2442 : inv port map( inb => mult_125_G3_ab_9_11_port, outb => n3955);
   U2443 : oai22 port map( a => n3953, b => n3955, c => n911, d => n2601, outb 
                           => n914);
   U2444 : aoi22 port map( a => n914, b => mult_125_G3_ab_10_11_port, c => 
                           n3957, d => n2604, outb => n3956);
   U2445 : inv port map( inb => mult_125_G3_ab_11_11_port, outb => n3958);
   U2446 : oai22 port map( a => n3956, b => n3958, c => n915, d => n2607, outb 
                           => n918);
   U2447 : aoi22 port map( a => n918, b => mult_125_G3_ab_12_11_port, c => 
                           n3960, d => n2610, outb => n3959);
   U2448 : inv port map( inb => mult_125_G3_ab_13_11_port, outb => n3961);
   U2449 : oai22 port map( a => n3959, b => n3961, c => n919, d => n2613, outb 
                           => n922);
   U2450 : aoi22 port map( a => n922, b => mult_125_G3_ab_14_11_port, c => 
                           n3962, d => n2616, outb => n925);
   U2451 : nand2 port map( a => mult_125_G3_ab_0_11_port, b => 
                           mult_125_G3_ab_1_10_port, outb => n928);
   U2452 : aoi22 port map( a => mult_125_G3_ab_2_10_port, b => n3964, c => n926
                           , d => n2584, outb => n3963);
   U2453 : oai22 port map( a => n3963, b => n3965, c => n929, d => n2585, outb 
                           => n932);
   U2454 : aoi22 port map( a => n932, b => mult_125_G3_ab_4_10_port, c => n3966
                           , d => n2624, outb => n935);
   U2455 : oai22 port map( a => n935, b => n934, c => n3967, d => n2587, outb 
                           => n937);
   U2456 : aoi22 port map( a => n937, b => mult_125_G3_ab_6_10_port, c => n3969
                           , d => n2627, outb => n3968);
   U2457 : oai22 port map( a => n3968, b => n3970, c => n938, d => n2590, outb 
                           => n941);
   U2458 : inv port map( inb => mult_125_G3_ab_8_10_port, outb => n3971);
   U2459 : oai22 port map( a => n3972, b => n3971, c => n940, d => n2593, outb 
                           => n943);
   U2460 : aoi22 port map( a => n943, b => mult_125_G3_ab_9_10_port, c => n3974
                           , d => n2596, outb => n3973);
   U2461 : inv port map( inb => mult_125_G3_ab_10_10_port, outb => n3975);
   U2462 : oai22 port map( a => n3973, b => n3975, c => n944, d => n2599, outb 
                           => n947);
   U2463 : aoi22 port map( a => n947, b => mult_125_G3_ab_11_10_port, c => 
                           n3977, d => n2602, outb => n3976);
   U2464 : inv port map( inb => mult_125_G3_ab_12_10_port, outb => n3978);
   U2465 : oai22 port map( a => n3976, b => n3978, c => n948, d => n2605, outb 
                           => n951);
   U2466 : aoi22 port map( a => n951, b => mult_125_G3_ab_13_10_port, c => 
                           n3980, d => n2608, outb => n3979);
   U2467 : inv port map( inb => mult_125_G3_ab_14_10_port, outb => n3981);
   U2468 : oai22 port map( a => n3979, b => n3981, c => n952, d => n2611, outb 
                           => n955);
   U2469 : nand2 port map( a => mult_125_G3_ab_0_10_port, b => 
                           mult_125_G3_ab_1_9_port, outb => n958);
   U2470 : aoi22 port map( a => mult_125_G3_ab_2_9_port, b => n3983, c => n956,
                           d => n2619, outb => n3982);
   U2471 : oai22 port map( a => n3982, b => n3984, c => n959, d => n2620, outb 
                           => n962);
   U2472 : oai22 port map( a => n3985, b => n3986, c => n961, d => n2633, outb 
                           => n964);
   U2473 : aoi22 port map( a => n964, b => mult_125_G3_ab_5_9_port, c => n3988,
                           d => n2622, outb => n3987);
   U2474 : oai22 port map( a => n3987, b => n3989, c => n965, d => n2636, outb 
                           => n968);
   U2475 : aoi22 port map( a => n968, b => mult_125_G3_ab_7_9_port, c => n3991,
                           d => n2625, outb => n3990);
   U2476 : oai22 port map( a => n3990, b => n3992, c => n969, d => n2639, outb 
                           => n972);
   U2477 : oai22 port map( a => n3993, b => n3994, c => n971, d => n2642, outb 
                           => n974);
   U2478 : aoi22 port map( a => n974, b => mult_125_G3_ab_10_9_port, c => n3996
                           , d => n2645, outb => n3995);
   U2479 : inv port map( inb => mult_125_G3_ab_11_9_port, outb => n3997);
   U2480 : oai22 port map( a => n3995, b => n3997, c => n975, d => n2648, outb 
                           => n978);
   U2481 : aoi22 port map( a => n978, b => mult_125_G3_ab_12_9_port, c => n3999
                           , d => n2651, outb => n3998);
   U2482 : inv port map( inb => mult_125_G3_ab_13_9_port, outb => n4000);
   U2483 : oai22 port map( a => n3998, b => n4000, c => n979, d => n2654, outb 
                           => n982);
   U2484 : aoi22 port map( a => n982, b => mult_125_G3_ab_14_9_port, c => n4001
                           , d => n2657, outb => n985);
   U2485 : nand2 port map( a => mult_125_G3_ab_0_9_port, b => 
                           mult_125_G3_ab_1_8_port, outb => n988);
   U2486 : aoi22 port map( a => mult_125_G3_ab_2_8_port, b => n4003, c => n986,
                           d => n2628, outb => n4002);
   U2487 : oai22 port map( a => n4002, b => n4004, c => n989, d => n2629, outb 
                           => n992);
   U2488 : oai22 port map( a => n4005, b => n4006, c => n991, d => n2665, outb 
                           => n994);
   U2489 : oai22 port map( a => n4007, b => n4008, c => n993, d => n2631, outb 
                           => n996);
   U2490 : aoi22 port map( a => n996, b => mult_125_G3_ab_6_8_port, c => n4010,
                           d => n2668, outb => n4009);
   U2491 : oai22 port map( a => n4009, b => n4011, c => n997, d => n2634, outb 
                           => n1000);
   U2492 : aoi22 port map( a => n1000, b => mult_125_G3_ab_8_8_port, c => n4013
                           , d => n2671, outb => n4012);
   U2493 : oai22 port map( a => n4012, b => n4014, c => n1001, d => n2637, outb
                           => n1004);
   U2494 : inv port map( inb => mult_125_G3_ab_10_8_port, outb => n4015);
   U2495 : oai22 port map( a => n4016, b => n4015, c => n1003, d => n2640, outb
                           => n1006);
   U2496 : aoi22 port map( a => n1006, b => mult_125_G3_ab_11_8_port, c => 
                           n4018, d => n2643, outb => n4017);
   U2497 : inv port map( inb => mult_125_G3_ab_12_8_port, outb => n4019);
   U2498 : oai22 port map( a => n4017, b => n4019, c => n1007, d => n2646, outb
                           => n1010);
   U2499 : aoi22 port map( a => n1010, b => mult_125_G3_ab_13_8_port, c => 
                           n4021, d => n2649, outb => n4020);
   U2500 : inv port map( inb => mult_125_G3_ab_14_8_port, outb => n4022);
   U2501 : oai22 port map( a => n4020, b => n4022, c => n1011, d => n2652, outb
                           => n1014);
   U2502 : nand2 port map( a => mult_125_G3_ab_0_8_port, b => 
                           mult_125_G3_ab_1_7_port, outb => n1017);
   U2503 : aoi22 port map( a => mult_125_G3_ab_2_7_port, b => n4023, c => n1015
                           , d => n2660, outb => n1020);
   U2504 : oai22 port map( a => n1020, b => n1019, c => n4024, d => n2661, outb
                           => n1022);
   U2505 : oai22 port map( a => n4025, b => n4026, c => n1021, d => n2677, outb
                           => n1024);
   U2506 : aoi22 port map( a => n1024, b => mult_125_G3_ab_5_7_port, c => n4028
                           , d => n2663, outb => n4027);
   U2507 : oai22 port map( a => n4027, b => n4029, c => n1025, d => n2680, outb
                           => n1028);
   U2508 : aoi22 port map( a => n1028, b => mult_125_G3_ab_7_7_port, c => n4031
                           , d => n2666, outb => n4030);
   U2509 : oai22 port map( a => n4030, b => n4032, c => n1029, d => n2683, outb
                           => n1032);
   U2510 : aoi22 port map( a => n1032, b => mult_125_G3_ab_9_7_port, c => n4034
                           , d => n2669, outb => n4033);
   U2511 : oai22 port map( a => n4033, b => n4035, c => n1033, d => n2686, outb
                           => n1036);
   U2512 : oai22 port map( a => n4036, b => n4037, c => n1035, d => n2689, outb
                           => n1038);
   U2513 : aoi22 port map( a => n1038, b => mult_125_G3_ab_12_7_port, c => 
                           n4039, d => n2692, outb => n4038);
   U2514 : inv port map( inb => mult_125_G3_ab_13_7_port, outb => n4040);
   U2515 : oai22 port map( a => n4038, b => n4040, c => n1039, d => n2695, outb
                           => n1042);
   U2516 : aoi22 port map( a => n1042, b => mult_125_G3_ab_14_7_port, c => 
                           n4041, d => n2698, outb => n1045);
   U2517 : nand2 port map( a => mult_125_G3_ab_0_7_port, b => 
                           mult_125_G3_ab_1_6_port, outb => n1048);
   U2518 : aoi22 port map( a => mult_125_G3_ab_2_6_port, b => n4043, c => n1046
                           , d => n2672, outb => n4042);
   U2519 : oai22 port map( a => n4042, b => n4044, c => n1049, d => n2673, outb
                           => n1052);
   U2520 : aoi22 port map( a => n1052, b => mult_125_G3_ab_4_6_port, c => n4045
                           , d => n2706, outb => n1055);
   U2521 : oai22 port map( a => n1055, b => n1054, c => n4046, d => n2675, outb
                           => n1057);
   U2522 : aoi22 port map( a => n1057, b => mult_125_G3_ab_6_6_port, c => n4048
                           , d => n2709, outb => n4047);
   U2523 : oai22 port map( a => n4047, b => n4049, c => n1058, d => n2678, outb
                           => n1061);
   U2524 : aoi22 port map( a => n1061, b => mult_125_G3_ab_8_6_port, c => n4050
                           , d => n2712, outb => n1064);
   U2525 : oai22 port map( a => n1064, b => n1063, c => n4051, d => n2681, outb
                           => n1066);
   U2526 : aoi22 port map( a => n1066, b => mult_125_G3_ab_10_6_port, c => 
                           n4053, d => n2715, outb => n4052);
   U2527 : oai22 port map( a => n4052, b => n4054, c => n1067, d => n2684, outb
                           => n1070);
   U2528 : inv port map( inb => mult_125_G3_ab_12_6_port, outb => n4055);
   U2529 : oai22 port map( a => n4056, b => n4055, c => n1069, d => n2687, outb
                           => n1072);
   U2530 : aoi22 port map( a => n1072, b => mult_125_G3_ab_13_6_port, c => 
                           n4058, d => n2690, outb => n4057);
   U2531 : inv port map( inb => mult_125_G3_ab_14_6_port, outb => n4059);
   U2532 : oai22 port map( a => n4057, b => n4059, c => n1073, d => n2693, outb
                           => n1076);
   U2533 : nand2 port map( a => mult_125_G3_ab_0_6_port, b => 
                           mult_125_G3_ab_1_5_port, outb => n1079);
   U2534 : aoi22 port map( a => mult_125_G3_ab_2_5_port, b => n4060, c => n1077
                           , d => n2701, outb => n1082);
   U2535 : oai22 port map( a => n1082, b => n1081, c => n4061, d => n2702, outb
                           => n1084);
   U2536 : oai22 port map( a => n4062, b => n4063, c => n1083, d => n2721, outb
                           => n1086);
   U2537 : aoi22 port map( a => n1086, b => mult_125_G3_ab_5_5_port, c => n4064
                           , d => n2704, outb => n1089);
   U2538 : oai22 port map( a => n1089, b => n1088, c => n4065, d => n2724, outb
                           => n1091);
   U2539 : aoi22 port map( a => n1091, b => mult_125_G3_ab_7_5_port, c => n4067
                           , d => n2707, outb => n4066);
   U2540 : oai22 port map( a => n4066, b => n4068, c => n1092, d => n2727, outb
                           => n1095);
   U2541 : aoi22 port map( a => n1095, b => mult_125_G3_ab_9_5_port, c => n4070
                           , d => n2710, outb => n4069);
   U2542 : oai22 port map( a => n4069, b => n4071, c => n1096, d => n2730, outb
                           => n1099);
   U2543 : aoi22 port map( a => n1099, b => mult_125_G3_ab_11_5_port, c => 
                           n4073, d => n2713, outb => n4072);
   U2544 : oai22 port map( a => n4072, b => n4074, c => n1100, d => n2733, outb
                           => n1103);
   U2545 : oai22 port map( a => n4075, b => n4076, c => n1102, d => n2736, outb
                           => n1105);
   U2546 : aoi22 port map( a => n1105, b => mult_125_G3_ab_14_5_port, c => 
                           n4077, d => n2739, outb => n1108);
   U2547 : nand2 port map( a => mult_125_G3_ab_0_5_port, b => 
                           mult_125_G3_ab_1_4_port, outb => n1111);
   U2548 : aoi22 port map( a => mult_125_G3_ab_2_4_port, b => n4079, c => n1109
                           , d => n2716, outb => n4078);
   U2549 : oai22 port map( a => n4078, b => n4080, c => n1112, d => n2717, outb
                           => n1115);
   U2550 : aoi22 port map( a => n1115, b => mult_125_G3_ab_4_4_port, c => n4081
                           , d => n2747, outb => n1118);
   U2551 : oai22 port map( a => n1118, b => n1117, c => n4082, d => n2719, outb
                           => n1120);
   U2552 : aoi22 port map( a => n1120, b => mult_125_G3_ab_6_4_port, c => n4083
                           , d => n2750, outb => n1123);
   U2553 : oai22 port map( a => n1123, b => n1122, c => n4084, d => n2722, outb
                           => n1125);
   U2554 : aoi22 port map( a => n1125, b => mult_125_G3_ab_8_4_port, c => n4086
                           , d => n2753, outb => n4085);
   U2555 : oai22 port map( a => n4085, b => n4087, c => n1126, d => n2725, outb
                           => n1129);
   U2556 : aoi22 port map( a => n1129, b => mult_125_G3_ab_10_4_port, c => 
                           n4088, d => n2756, outb => n1132);
   U2557 : oai22 port map( a => n1132, b => n1131, c => n4089, d => n2728, outb
                           => n1134);
   U2558 : aoi22 port map( a => n1134, b => mult_125_G3_ab_12_4_port, c => 
                           n4091, d => n2759, outb => n4090);
   U2559 : oai22 port map( a => n4090, b => n4092, c => n1135, d => n2731, outb
                           => n1138);
   U2560 : aoi22 port map( a => n1138, b => mult_125_G3_ab_14_4_port, c => 
                           n4093, d => n2734, outb => n1141);
   U2561 : nand2 port map( a => mult_125_G3_ab_0_4_port, b => 
                           mult_125_G3_ab_1_3_port, outb => n1144);
   U2562 : aoi22 port map( a => mult_125_G3_ab_2_3_port, b => n4094, c => n1142
                           , d => n2742, outb => n1147);
   U2563 : oai22 port map( a => n1147, b => n1146, c => n4095, d => n2743, outb
                           => n1149);
   U2564 : oai22 port map( a => n4096, b => n4097, c => n1148, d => n2765, outb
                           => n1151);
   U2565 : aoi22 port map( a => n1151, b => mult_125_G3_ab_5_3_port, c => n4099
                           , d => n2745, outb => n4098);
   U2566 : oai22 port map( a => n4098, b => n4100, c => n1152, d => n2768, outb
                           => n1155);
   U2567 : aoi22 port map( a => n1155, b => mult_125_G3_ab_7_3_port, c => n4102
                           , d => n2748, outb => n4101);
   U2568 : oai22 port map( a => n4101, b => n4103, c => n1156, d => n2771, outb
                           => n1159);
   U2569 : aoi22 port map( a => n1159, b => mult_125_G3_ab_9_3_port, c => n4105
                           , d => n2751, outb => n4104);
   U2570 : oai22 port map( a => n4104, b => n4106, c => n1160, d => n2774, outb
                           => n1163);
   U2571 : aoi22 port map( a => n1163, b => mult_125_G3_ab_11_3_port, c => 
                           n4108, d => n2754, outb => n4107);
   U2572 : oai22 port map( a => n4107, b => n4109, c => n1164, d => n2777, outb
                           => n1167);
   U2573 : aoi22 port map( a => n1167, b => mult_125_G3_ab_13_3_port, c => 
                           n4111, d => n2757, outb => n4110);
   U2574 : inv port map( inb => mult_125_G3_ab_14_3_port, outb => n4112);
   U2575 : oai22 port map( a => n4110, b => n4112, c => n1168, d => n2780, outb
                           => n1171);
   U2576 : nand2 port map( a => mult_125_G3_ab_0_3_port, b => 
                           mult_125_G3_ab_1_2_port, outb => n1174);
   U2577 : aoi22 port map( a => mult_125_G3_ab_2_2_port, b => n4114, c => n1172
                           , d => n2760, outb => n4113);
   U2578 : oai22 port map( a => n4113, b => n4115, c => n1175, d => n2761, outb
                           => n1178);
   U2579 : aoi22 port map( a => n1178, b => mult_125_G3_ab_4_2_port, c => n4117
                           , d => n2788, outb => n4116);
   U2580 : oai22 port map( a => n4116, b => n4118, c => n1179, d => n2763, outb
                           => n1182);
   U2581 : aoi22 port map( a => n1182, b => mult_125_G3_ab_6_2_port, c => n4119
                           , d => n2791, outb => n1185);
   U2582 : oai22 port map( a => n1185, b => n1184, c => n4120, d => n2766, outb
                           => n1187);
   U2583 : aoi22 port map( a => n1187, b => mult_125_G3_ab_8_2_port, c => n4122
                           , d => n2794, outb => n4121);
   U2584 : oai22 port map( a => n4121, b => n4123, c => n1188, d => n2769, outb
                           => n1191);
   U2585 : aoi22 port map( a => n1191, b => mult_125_G3_ab_10_2_port, c => 
                           n4125, d => n2797, outb => n4124);
   U2586 : oai22 port map( a => n4124, b => n4126, c => n1192, d => n2772, outb
                           => n1195);
   U2587 : aoi22 port map( a => n1195, b => mult_125_G3_ab_12_2_port, c => 
                           n4128, d => n2800, outb => n4127);
   U2588 : oai22 port map( a => n4127, b => n4129, c => n1196, d => n2775, outb
                           => n1199);
   U2589 : aoi22 port map( a => n1199, b => mult_125_G3_ab_14_2_port, c => 
                           n4131, d => n2803, outb => n4130);
   U2590 : nand2 port map( a => mult_125_G3_ab_0_2_port, b => 
                           mult_125_G3_ab_1_1_port, outb => n1204);
   U2591 : aoi22 port map( a => mult_125_G3_ab_2_1_port, b => n4133, c => n1202
                           , d => n2783, outb => n4132);
   U2592 : oai22 port map( a => n4132, b => n4134, c => n1205, d => n2784, outb
                           => n1208);
   U2593 : inv port map( inb => mult_125_G3_ab_4_1_port, outb => n4135);
   U2594 : oai22 port map( a => n4136, b => n4135, c => n1207, d => n2809, outb
                           => n1210);
   U2595 : aoi22 port map( a => n1210, b => mult_125_G3_ab_5_1_port, c => n4138
                           , d => n2786, outb => n4137);
   U2596 : oai22 port map( a => n4137, b => n4139, c => n1211, d => n2812, outb
                           => n1214);
   U2597 : aoi22 port map( a => n1214, b => mult_125_G3_ab_7_1_port, c => n4141
                           , d => n2789, outb => n4140);
   U2598 : oai22 port map( a => n4140, b => n4142, c => n1215, d => n2815, outb
                           => n1218);
   U2599 : aoi22 port map( a => n1218, b => mult_125_G3_ab_9_1_port, c => n4144
                           , d => n2792, outb => n4143);
   U2600 : oai22 port map( a => n4143, b => n4145, c => n1219, d => n2818, outb
                           => n1222);
   U2601 : aoi22 port map( a => n1222, b => mult_125_G3_ab_11_1_port, c => 
                           n4147, d => n2795, outb => n4146);
   U2602 : oai22 port map( a => n4146, b => n4148, c => n1223, d => n2821, outb
                           => n1226);
   U2603 : aoi22 port map( a => n1226, b => mult_125_G3_ab_13_1_port, c => 
                           n4150, d => n2798, outb => n4149);
   U2604 : inv port map( inb => mult_125_G3_ab_14_1_port, outb => n4151);
   U2605 : oai22 port map( a => n4149, b => n4151, c => n1227, d => n2824, outb
                           => n1230);
   U2606 : nand2 port map( a => mult_125_G3_ab_0_1_port, b => 
                           mult_125_G3_ab_1_0_port, outb => n4152);
   U2607 : aoi22 port map( a => mult_125_G3_ab_2_0_port, b => n1232, c => n4154
                           , d => n2804, outb => n4153);
   U2608 : aoi22 port map( a => n1234, b => mult_125_G3_ab_3_0_port, c => n4156
                           , d => n2805, outb => n4155);
   U2609 : inv port map( inb => mult_125_G3_ab_4_0_port, outb => n4157);
   U2610 : oai22 port map( a => n4155, b => n4157, c => n1235, d => n4158, outb
                           => n1238);
   U2611 : aoi22 port map( a => n1238, b => mult_125_G3_ab_5_0_port, c => n4160
                           , d => n2807, outb => n4159);
   U2612 : inv port map( inb => mult_125_G3_ab_6_0_port, outb => n4161);
   U2613 : oai22 port map( a => n4159, b => n4161, c => n1239, d => n4162, outb
                           => n1242);
   U2614 : aoi22 port map( a => n1242, b => mult_125_G3_ab_7_0_port, c => n4164
                           , d => n2810, outb => n4163);
   U2615 : inv port map( inb => mult_125_G3_ab_8_0_port, outb => n4165);
   U2616 : oai22 port map( a => n4163, b => n4165, c => n1243, d => n4166, outb
                           => n1246);
   U2617 : aoi22 port map( a => n1246, b => mult_125_G3_ab_9_0_port, c => n4168
                           , d => n2813, outb => n4167);
   U2618 : inv port map( inb => mult_125_G3_ab_10_0_port, outb => n4169);
   U2619 : oai22 port map( a => n4167, b => n4169, c => n1247, d => n4170, outb
                           => n1250);
   U2620 : aoi22 port map( a => n1250, b => mult_125_G3_ab_11_0_port, c => 
                           n4172, d => n2816, outb => n4171);
   U2621 : inv port map( inb => mult_125_G3_ab_12_0_port, outb => n4173);
   U2622 : oai22 port map( a => n4171, b => n4173, c => n1251, d => n4174, outb
                           => n1254);
   U2623 : aoi22 port map( a => n1254, b => mult_125_G3_ab_13_0_port, c => 
                           n4176, d => n2819, outb => n4175);
   U2624 : inv port map( inb => mult_125_G3_ab_14_0_port, outb => n4177);
   U2625 : oai22 port map( a => n4175, b => n4177, c => n1255, d => n4178, outb
                           => n1258);
   U2626 : inv port map( inb => mult_125_G3_ZB, outb => n380);
   U2627 : inv port map( inb => mult_125_G3_ZA, outb => n381);
   U2628 : nand2 port map( a => mult_125_G2_ab_0_15_port, b => 
                           mult_125_G2_ab_1_14_port, outb => n4179);
   U2629 : inv port map( inb => mult_125_G2_ab_3_15_port, outb => n4180);
   U2630 : inv port map( inb => mult_125_G2_ab_4_14_port, outb => n4181);
   U2631 : inv port map( inb => mult_125_G2_ab_5_15_port, outb => n4182);
   U2632 : inv port map( inb => mult_125_G2_ab_6_14_port, outb => n4183);
   U2633 : inv port map( inb => mult_125_G2_ab_7_15_port, outb => n4184);
   U2634 : inv port map( inb => mult_125_G2_ab_8_14_port, outb => n4185);
   U2635 : inv port map( inb => mult_125_G2_ab_9_15_port, outb => n4186);
   U2636 : inv port map( inb => mult_125_G2_ab_10_14_port, outb => n4187);
   U2637 : inv port map( inb => mult_125_G2_ab_11_15_port, outb => n4188);
   U2638 : inv port map( inb => mult_125_G2_ab_12_14_port, outb => n4189);
   U2639 : nand2 port map( a => mult_125_G2_ab_0_14_port, b => 
                           mult_125_G2_ab_1_13_port, outb => n1276);
   U2640 : aoi22 port map( a => mult_125_G2_ab_2_13_port, b => n4190, c => 
                           n1274, d => n2834, outb => n1279);
   U2641 : oai22 port map( a => n1279, b => n1278, c => n4191, d => n2835, outb
                           => n1281);
   U2642 : aoi22 port map( a => n1281, b => mult_125_G2_ab_4_13_port, c => 
                           n4193, d => n2842, outb => n4192);
   U2643 : oai22 port map( a => n4192, b => n4194, c => n1282, d => n2845, outb
                           => n1285);
   U2644 : aoi22 port map( a => n1285, b => mult_125_G2_ab_6_13_port, c => 
                           n4196, d => n2848, outb => n4195);
   U2645 : inv port map( inb => mult_125_G2_ab_7_13_port, outb => n4197);
   U2646 : oai22 port map( a => n4195, b => n4197, c => n1286, d => n2851, outb
                           => n1289);
   U2647 : aoi22 port map( a => n1289, b => mult_125_G2_ab_8_13_port, c => 
                           n4199, d => n2854, outb => n4198);
   U2648 : inv port map( inb => mult_125_G2_ab_9_13_port, outb => n4200);
   U2649 : oai22 port map( a => n4198, b => n4200, c => n1290, d => n2857, outb
                           => n1293);
   U2650 : aoi22 port map( a => n1293, b => mult_125_G2_ab_10_13_port, c => 
                           n4202, d => n2860, outb => n4201);
   U2651 : inv port map( inb => mult_125_G2_ab_11_13_port, outb => n4203);
   U2652 : oai22 port map( a => n4201, b => n4203, c => n1294, d => n2863, outb
                           => n1297);
   U2653 : aoi22 port map( a => n1297, b => mult_125_G2_ab_12_13_port, c => 
                           n4205, d => n2866, outb => n4204);
   U2654 : inv port map( inb => mult_125_G2_ab_13_13_port, outb => n4206);
   U2655 : oai22 port map( a => n4204, b => n4206, c => n1298, d => n2869, outb
                           => n1301);
   U2656 : aoi22 port map( a => n1301, b => mult_125_G2_ab_14_13_port, c => 
                           n4208, d => n2872, outb => n4207);
   U2657 : nand2 port map( a => mult_125_G2_ab_0_13_port, b => 
                           mult_125_G2_ab_1_12_port, outb => n1306);
   U2658 : aoi22 port map( a => mult_125_G2_ab_2_12_port, b => n4210, c => 
                           n1304, d => n2837, outb => n4209);
   U2659 : oai22 port map( a => n4209, b => n4211, c => n1307, d => n2838, outb
                           => n1310);
   U2660 : aoi22 port map( a => n1310, b => mult_125_G2_ab_4_12_port, c => 
                           n4213, d => n2880, outb => n4212);
   U2661 : aoi22 port map( a => n1312, b => mult_125_G2_ab_5_12_port, c => 
                           n4215, d => n2840, outb => n4214);
   U2662 : inv port map( inb => mult_125_G2_ab_6_12_port, outb => n4216);
   U2663 : oai22 port map( a => n4214, b => n4216, c => n1313, d => n2843, outb
                           => n1316);
   U2664 : aoi22 port map( a => n1316, b => mult_125_G2_ab_7_12_port, c => 
                           n4218, d => n2846, outb => n4217);
   U2665 : inv port map( inb => mult_125_G2_ab_8_12_port, outb => n4219);
   U2666 : oai22 port map( a => n4217, b => n4219, c => n1317, d => n2849, outb
                           => n1320);
   U2667 : aoi22 port map( a => n1320, b => mult_125_G2_ab_9_12_port, c => 
                           n4221, d => n2852, outb => n4220);
   U2668 : inv port map( inb => mult_125_G2_ab_10_12_port, outb => n4222);
   U2669 : oai22 port map( a => n4220, b => n4222, c => n1321, d => n2855, outb
                           => n1324);
   U2670 : aoi22 port map( a => n1324, b => mult_125_G2_ab_11_12_port, c => 
                           n4224, d => n2858, outb => n4223);
   U2671 : inv port map( inb => mult_125_G2_ab_12_12_port, outb => n4225);
   U2672 : oai22 port map( a => n4223, b => n4225, c => n1325, d => n2861, outb
                           => n1328);
   U2673 : aoi22 port map( a => n1328, b => mult_125_G2_ab_13_12_port, c => 
                           n4227, d => n2864, outb => n4226);
   U2674 : inv port map( inb => mult_125_G2_ab_14_12_port, outb => n4228);
   U2675 : oai22 port map( a => n4226, b => n4228, c => n1329, d => n2867, outb
                           => n1332);
   U2676 : nand2 port map( a => mult_125_G2_ab_0_12_port, b => 
                           mult_125_G2_ab_1_11_port, outb => n1335);
   U2677 : aoi22 port map( a => mult_125_G2_ab_2_11_port, b => n4229, c => 
                           n1333, d => n2875, outb => n1338);
   U2678 : oai22 port map( a => n1338, b => n1337, c => n4230, d => n2876, outb
                           => n1340);
   U2679 : oai22 port map( a => n4231, b => n4232, c => n1339, d => n2886, outb
                           => n1342);
   U2680 : aoi22 port map( a => n1342, b => mult_125_G2_ab_5_11_port, c => 
                           n4234, d => n2878, outb => n4233);
   U2681 : oai22 port map( a => n4233, b => n4235, c => n1343, d => n2889, outb
                           => n1346);
   U2682 : oai22 port map( a => n4236, b => n4237, c => n1345, d => n2892, outb
                           => n1348);
   U2683 : aoi22 port map( a => n1348, b => mult_125_G2_ab_8_11_port, c => 
                           n4239, d => n2895, outb => n4238);
   U2684 : inv port map( inb => mult_125_G2_ab_9_11_port, outb => n4240);
   U2685 : oai22 port map( a => n4238, b => n4240, c => n1349, d => n2898, outb
                           => n1352);
   U2686 : aoi22 port map( a => n1352, b => mult_125_G2_ab_10_11_port, c => 
                           n4242, d => n2901, outb => n4241);
   U2687 : inv port map( inb => mult_125_G2_ab_11_11_port, outb => n4243);
   U2688 : oai22 port map( a => n4241, b => n4243, c => n1353, d => n2904, outb
                           => n1356);
   U2689 : aoi22 port map( a => n1356, b => mult_125_G2_ab_12_11_port, c => 
                           n4245, d => n2907, outb => n4244);
   U2690 : inv port map( inb => mult_125_G2_ab_13_11_port, outb => n4246);
   U2691 : oai22 port map( a => n4244, b => n4246, c => n1357, d => n2910, outb
                           => n1360);
   U2692 : aoi22 port map( a => n1360, b => mult_125_G2_ab_14_11_port, c => 
                           n4247, d => n2913, outb => n1363);
   U2693 : nand2 port map( a => mult_125_G2_ab_0_11_port, b => 
                           mult_125_G2_ab_1_10_port, outb => n1366);
   U2694 : aoi22 port map( a => mult_125_G2_ab_2_10_port, b => n4249, c => 
                           n1364, d => n2881, outb => n4248);
   U2695 : oai22 port map( a => n4248, b => n4250, c => n1367, d => n2882, outb
                           => n1370);
   U2696 : aoi22 port map( a => n1370, b => mult_125_G2_ab_4_10_port, c => 
                           n4251, d => n2921, outb => n1373);
   U2697 : oai22 port map( a => n1373, b => n1372, c => n4252, d => n2884, outb
                           => n1375);
   U2698 : aoi22 port map( a => n1375, b => mult_125_G2_ab_6_10_port, c => 
                           n4254, d => n2924, outb => n4253);
   U2699 : oai22 port map( a => n4253, b => n4255, c => n1376, d => n2887, outb
                           => n1379);
   U2700 : inv port map( inb => mult_125_G2_ab_8_10_port, outb => n4256);
   U2701 : oai22 port map( a => n4257, b => n4256, c => n1378, d => n2890, outb
                           => n1381);
   U2702 : aoi22 port map( a => n1381, b => mult_125_G2_ab_9_10_port, c => 
                           n4259, d => n2893, outb => n4258);
   U2703 : inv port map( inb => mult_125_G2_ab_10_10_port, outb => n4260);
   U2704 : oai22 port map( a => n4258, b => n4260, c => n1382, d => n2896, outb
                           => n1385);
   U2705 : aoi22 port map( a => n1385, b => mult_125_G2_ab_11_10_port, c => 
                           n4262, d => n2899, outb => n4261);
   U2706 : inv port map( inb => mult_125_G2_ab_12_10_port, outb => n4263);
   U2707 : oai22 port map( a => n4261, b => n4263, c => n1386, d => n2902, outb
                           => n1389);
   U2708 : aoi22 port map( a => n1389, b => mult_125_G2_ab_13_10_port, c => 
                           n4265, d => n2905, outb => n4264);
   U2709 : inv port map( inb => mult_125_G2_ab_14_10_port, outb => n4266);
   U2710 : oai22 port map( a => n4264, b => n4266, c => n1390, d => n2908, outb
                           => n1393);
   U2711 : nand2 port map( a => mult_125_G2_ab_0_10_port, b => 
                           mult_125_G2_ab_1_9_port, outb => n1396);
   U2712 : aoi22 port map( a => mult_125_G2_ab_2_9_port, b => n4268, c => n1394
                           , d => n2916, outb => n4267);
   U2713 : oai22 port map( a => n4267, b => n4269, c => n1397, d => n2917, outb
                           => n1400);
   U2714 : oai22 port map( a => n4270, b => n4271, c => n1399, d => n2930, outb
                           => n1402);
   U2715 : aoi22 port map( a => n1402, b => mult_125_G2_ab_5_9_port, c => n4273
                           , d => n2919, outb => n4272);
   U2716 : oai22 port map( a => n4272, b => n4274, c => n1403, d => n2933, outb
                           => n1406);
   U2717 : aoi22 port map( a => n1406, b => mult_125_G2_ab_7_9_port, c => n4276
                           , d => n2922, outb => n4275);
   U2718 : oai22 port map( a => n4275, b => n4277, c => n1407, d => n2936, outb
                           => n1410);
   U2719 : oai22 port map( a => n4278, b => n4279, c => n1409, d => n2939, outb
                           => n1412);
   U2720 : aoi22 port map( a => n1412, b => mult_125_G2_ab_10_9_port, c => 
                           n4281, d => n2942, outb => n4280);
   U2721 : inv port map( inb => mult_125_G2_ab_11_9_port, outb => n4282);
   U2722 : oai22 port map( a => n4280, b => n4282, c => n1413, d => n2945, outb
                           => n1416);
   U2723 : aoi22 port map( a => n1416, b => mult_125_G2_ab_12_9_port, c => 
                           n4284, d => n2948, outb => n4283);
   U2724 : inv port map( inb => mult_125_G2_ab_13_9_port, outb => n4285);
   U2725 : oai22 port map( a => n4283, b => n4285, c => n1417, d => n2951, outb
                           => n1420);
   U2726 : aoi22 port map( a => n1420, b => mult_125_G2_ab_14_9_port, c => 
                           n4286, d => n2954, outb => n1423);
   U2727 : nand2 port map( a => mult_125_G2_ab_0_9_port, b => 
                           mult_125_G2_ab_1_8_port, outb => n1426);
   U2728 : aoi22 port map( a => mult_125_G2_ab_2_8_port, b => n4288, c => n1424
                           , d => n2925, outb => n4287);
   U2729 : oai22 port map( a => n4287, b => n4289, c => n1427, d => n2926, outb
                           => n1430);
   U2730 : oai22 port map( a => n4290, b => n4291, c => n1429, d => n2962, outb
                           => n1432);
   U2731 : oai22 port map( a => n4292, b => n4293, c => n1431, d => n2928, outb
                           => n1434);
   U2732 : aoi22 port map( a => n1434, b => mult_125_G2_ab_6_8_port, c => n4295
                           , d => n2965, outb => n4294);
   U2733 : oai22 port map( a => n4294, b => n4296, c => n1435, d => n2931, outb
                           => n1438);
   U2734 : aoi22 port map( a => n1438, b => mult_125_G2_ab_8_8_port, c => n4298
                           , d => n2968, outb => n4297);
   U2735 : oai22 port map( a => n4297, b => n4299, c => n1439, d => n2934, outb
                           => n1442);
   U2736 : inv port map( inb => mult_125_G2_ab_10_8_port, outb => n4300);
   U2737 : oai22 port map( a => n4301, b => n4300, c => n1441, d => n2937, outb
                           => n1444);
   U2738 : aoi22 port map( a => n1444, b => mult_125_G2_ab_11_8_port, c => 
                           n4303, d => n2940, outb => n4302);
   U2739 : inv port map( inb => mult_125_G2_ab_12_8_port, outb => n4304);
   U2740 : oai22 port map( a => n4302, b => n4304, c => n1445, d => n2943, outb
                           => n1448);
   U2741 : aoi22 port map( a => n1448, b => mult_125_G2_ab_13_8_port, c => 
                           n4306, d => n2946, outb => n4305);
   U2742 : inv port map( inb => mult_125_G2_ab_14_8_port, outb => n4307);
   U2743 : oai22 port map( a => n4305, b => n4307, c => n1449, d => n2949, outb
                           => n1452);
   U2744 : nand2 port map( a => mult_125_G2_ab_0_8_port, b => 
                           mult_125_G2_ab_1_7_port, outb => n1455);
   U2745 : aoi22 port map( a => mult_125_G2_ab_2_7_port, b => n4308, c => n1453
                           , d => n2957, outb => n1458);
   U2746 : oai22 port map( a => n1458, b => n1457, c => n4309, d => n2958, outb
                           => n1460);
   U2747 : oai22 port map( a => n4310, b => n4311, c => n1459, d => n2974, outb
                           => n1462);
   U2748 : aoi22 port map( a => n1462, b => mult_125_G2_ab_5_7_port, c => n4313
                           , d => n2960, outb => n4312);
   U2749 : oai22 port map( a => n4312, b => n4314, c => n1463, d => n2977, outb
                           => n1466);
   U2750 : aoi22 port map( a => n1466, b => mult_125_G2_ab_7_7_port, c => n4316
                           , d => n2963, outb => n4315);
   U2751 : oai22 port map( a => n4315, b => n4317, c => n1467, d => n2980, outb
                           => n1470);
   U2752 : aoi22 port map( a => n1470, b => mult_125_G2_ab_9_7_port, c => n4319
                           , d => n2966, outb => n4318);
   U2753 : oai22 port map( a => n4318, b => n4320, c => n1471, d => n2983, outb
                           => n1474);
   U2754 : oai22 port map( a => n4321, b => n4322, c => n1473, d => n2986, outb
                           => n1476);
   U2755 : aoi22 port map( a => n1476, b => mult_125_G2_ab_12_7_port, c => 
                           n4324, d => n2989, outb => n4323);
   U2756 : inv port map( inb => mult_125_G2_ab_13_7_port, outb => n4325);
   U2757 : oai22 port map( a => n4323, b => n4325, c => n1477, d => n2992, outb
                           => n1480);
   U2758 : aoi22 port map( a => n1480, b => mult_125_G2_ab_14_7_port, c => 
                           n4326, d => n2995, outb => n1483);
   U2759 : nand2 port map( a => mult_125_G2_ab_0_7_port, b => 
                           mult_125_G2_ab_1_6_port, outb => n1486);
   U2760 : aoi22 port map( a => mult_125_G2_ab_2_6_port, b => n4328, c => n1484
                           , d => n2969, outb => n4327);
   U2761 : oai22 port map( a => n4327, b => n4329, c => n1487, d => n2970, outb
                           => n1490);
   U2762 : aoi22 port map( a => n1490, b => mult_125_G2_ab_4_6_port, c => n4330
                           , d => n3003, outb => n1493);
   U2763 : oai22 port map( a => n1493, b => n1492, c => n4331, d => n2972, outb
                           => n1495);
   U2764 : aoi22 port map( a => n1495, b => mult_125_G2_ab_6_6_port, c => n4333
                           , d => n3006, outb => n4332);
   U2765 : oai22 port map( a => n4332, b => n4334, c => n1496, d => n2975, outb
                           => n1499);
   U2766 : aoi22 port map( a => n1499, b => mult_125_G2_ab_8_6_port, c => n4335
                           , d => n3009, outb => n1502);
   U2767 : oai22 port map( a => n1502, b => n1501, c => n4336, d => n2978, outb
                           => n1504);
   U2768 : aoi22 port map( a => n1504, b => mult_125_G2_ab_10_6_port, c => 
                           n4338, d => n3012, outb => n4337);
   U2769 : oai22 port map( a => n4337, b => n4339, c => n1505, d => n2981, outb
                           => n1508);
   U2770 : inv port map( inb => mult_125_G2_ab_12_6_port, outb => n4340);
   U2771 : oai22 port map( a => n4341, b => n4340, c => n1507, d => n2984, outb
                           => n1510);
   U2772 : aoi22 port map( a => n1510, b => mult_125_G2_ab_13_6_port, c => 
                           n4343, d => n2987, outb => n4342);
   U2773 : inv port map( inb => mult_125_G2_ab_14_6_port, outb => n4344);
   U2774 : oai22 port map( a => n4342, b => n4344, c => n1511, d => n2990, outb
                           => n1514);
   U2775 : nand2 port map( a => mult_125_G2_ab_0_6_port, b => 
                           mult_125_G2_ab_1_5_port, outb => n1517);
   U2776 : aoi22 port map( a => mult_125_G2_ab_2_5_port, b => n4345, c => n1515
                           , d => n2998, outb => n1520);
   U2777 : oai22 port map( a => n1520, b => n1519, c => n4346, d => n2999, outb
                           => n1522);
   U2778 : oai22 port map( a => n4347, b => n4348, c => n1521, d => n3018, outb
                           => n1524);
   U2779 : aoi22 port map( a => n1524, b => mult_125_G2_ab_5_5_port, c => n4349
                           , d => n3001, outb => n1527);
   U2780 : oai22 port map( a => n1527, b => n1526, c => n4350, d => n3021, outb
                           => n1529);
   U2781 : aoi22 port map( a => n1529, b => mult_125_G2_ab_7_5_port, c => n4352
                           , d => n3004, outb => n4351);
   U2782 : oai22 port map( a => n4351, b => n4353, c => n1530, d => n3024, outb
                           => n1533);
   U2783 : aoi22 port map( a => n1533, b => mult_125_G2_ab_9_5_port, c => n4355
                           , d => n3007, outb => n4354);
   U2784 : oai22 port map( a => n4354, b => n4356, c => n1534, d => n3027, outb
                           => n1537);
   U2785 : aoi22 port map( a => n1537, b => mult_125_G2_ab_11_5_port, c => 
                           n4358, d => n3010, outb => n4357);
   U2786 : oai22 port map( a => n4357, b => n4359, c => n1538, d => n3030, outb
                           => n1541);
   U2787 : oai22 port map( a => n4360, b => n4361, c => n1540, d => n3033, outb
                           => n1543);
   U2788 : aoi22 port map( a => n1543, b => mult_125_G2_ab_14_5_port, c => 
                           n4362, d => n3036, outb => n1546);
   U2789 : nand2 port map( a => mult_125_G2_ab_0_5_port, b => 
                           mult_125_G2_ab_1_4_port, outb => n1549);
   U2790 : aoi22 port map( a => mult_125_G2_ab_2_4_port, b => n4364, c => n1547
                           , d => n3013, outb => n4363);
   U2791 : oai22 port map( a => n4363, b => n4365, c => n1550, d => n3014, outb
                           => n1553);
   U2792 : aoi22 port map( a => n1553, b => mult_125_G2_ab_4_4_port, c => n4366
                           , d => n3044, outb => n1556);
   U2793 : oai22 port map( a => n1556, b => n1555, c => n4367, d => n3016, outb
                           => n1558);
   U2794 : aoi22 port map( a => n1558, b => mult_125_G2_ab_6_4_port, c => n4368
                           , d => n3047, outb => n1561);
   U2795 : oai22 port map( a => n1561, b => n1560, c => n4369, d => n3019, outb
                           => n1563);
   U2796 : aoi22 port map( a => n1563, b => mult_125_G2_ab_8_4_port, c => n4371
                           , d => n3050, outb => n4370);
   U2797 : oai22 port map( a => n4370, b => n4372, c => n1564, d => n3022, outb
                           => n1567);
   U2798 : aoi22 port map( a => n1567, b => mult_125_G2_ab_10_4_port, c => 
                           n4373, d => n3053, outb => n1570);
   U2799 : oai22 port map( a => n1570, b => n1569, c => n4374, d => n3025, outb
                           => n1572);
   U2800 : aoi22 port map( a => n1572, b => mult_125_G2_ab_12_4_port, c => 
                           n4376, d => n3056, outb => n4375);
   U2801 : oai22 port map( a => n4375, b => n4377, c => n1573, d => n3028, outb
                           => n1576);
   U2802 : aoi22 port map( a => n1576, b => mult_125_G2_ab_14_4_port, c => 
                           n4378, d => n3031, outb => n1579);
   U2803 : nand2 port map( a => mult_125_G2_ab_0_4_port, b => 
                           mult_125_G2_ab_1_3_port, outb => n1582);
   U2804 : aoi22 port map( a => mult_125_G2_ab_2_3_port, b => n4379, c => n1580
                           , d => n3039, outb => n1585);
   U2805 : oai22 port map( a => n1585, b => n1584, c => n4380, d => n3040, outb
                           => n1587);
   U2806 : oai22 port map( a => n4381, b => n4382, c => n1586, d => n3062, outb
                           => n1589);
   U2807 : aoi22 port map( a => n1589, b => mult_125_G2_ab_5_3_port, c => n4384
                           , d => n3042, outb => n4383);
   U2808 : oai22 port map( a => n4383, b => n4385, c => n1590, d => n3065, outb
                           => n1593);
   U2809 : aoi22 port map( a => n1593, b => mult_125_G2_ab_7_3_port, c => n4387
                           , d => n3045, outb => n4386);
   U2810 : oai22 port map( a => n4386, b => n4388, c => n1594, d => n3068, outb
                           => n1597);
   U2811 : aoi22 port map( a => n1597, b => mult_125_G2_ab_9_3_port, c => n4390
                           , d => n3048, outb => n4389);
   U2812 : oai22 port map( a => n4389, b => n4391, c => n1598, d => n3071, outb
                           => n1601);
   U2813 : aoi22 port map( a => n1601, b => mult_125_G2_ab_11_3_port, c => 
                           n4393, d => n3051, outb => n4392);
   U2814 : oai22 port map( a => n4392, b => n4394, c => n1602, d => n3074, outb
                           => n1605);
   U2815 : aoi22 port map( a => n1605, b => mult_125_G2_ab_13_3_port, c => 
                           n4396, d => n3054, outb => n4395);
   U2816 : inv port map( inb => mult_125_G2_ab_14_3_port, outb => n4397);
   U2817 : oai22 port map( a => n4395, b => n4397, c => n1606, d => n3077, outb
                           => n1609);
   U2818 : nand2 port map( a => mult_125_G2_ab_0_3_port, b => 
                           mult_125_G2_ab_1_2_port, outb => n1612);
   U2819 : aoi22 port map( a => mult_125_G2_ab_2_2_port, b => n4399, c => n1610
                           , d => n3057, outb => n4398);
   U2820 : oai22 port map( a => n4398, b => n4400, c => n1613, d => n3058, outb
                           => n1616);
   U2821 : aoi22 port map( a => n1616, b => mult_125_G2_ab_4_2_port, c => n4402
                           , d => n3085, outb => n4401);
   U2822 : oai22 port map( a => n4401, b => n4403, c => n1617, d => n3060, outb
                           => n1620);
   U2823 : aoi22 port map( a => n1620, b => mult_125_G2_ab_6_2_port, c => n4404
                           , d => n3088, outb => n1623);
   U2824 : oai22 port map( a => n1623, b => n1622, c => n4405, d => n3063, outb
                           => n1625);
   U2825 : aoi22 port map( a => n1625, b => mult_125_G2_ab_8_2_port, c => n4407
                           , d => n3091, outb => n4406);
   U2826 : oai22 port map( a => n4406, b => n4408, c => n1626, d => n3066, outb
                           => n1629);
   U2827 : aoi22 port map( a => n1629, b => mult_125_G2_ab_10_2_port, c => 
                           n4410, d => n3094, outb => n4409);
   U2828 : oai22 port map( a => n4409, b => n4411, c => n1630, d => n3069, outb
                           => n1633);
   U2829 : aoi22 port map( a => n1633, b => mult_125_G2_ab_12_2_port, c => 
                           n4413, d => n3097, outb => n4412);
   U2830 : oai22 port map( a => n4412, b => n4414, c => n1634, d => n3072, outb
                           => n1637);
   U2831 : aoi22 port map( a => n1637, b => mult_125_G2_ab_14_2_port, c => 
                           n4416, d => n3100, outb => n4415);
   U2832 : nand2 port map( a => mult_125_G2_ab_0_2_port, b => 
                           mult_125_G2_ab_1_1_port, outb => n1642);
   U2833 : aoi22 port map( a => mult_125_G2_ab_2_1_port, b => n4418, c => n1640
                           , d => n3080, outb => n4417);
   U2834 : oai22 port map( a => n4417, b => n4419, c => n1643, d => n3081, outb
                           => n1646);
   U2835 : inv port map( inb => mult_125_G2_ab_4_1_port, outb => n4420);
   U2836 : oai22 port map( a => n4421, b => n4420, c => n1645, d => n3106, outb
                           => n1648);
   U2837 : aoi22 port map( a => n1648, b => mult_125_G2_ab_5_1_port, c => n4423
                           , d => n3083, outb => n4422);
   U2838 : oai22 port map( a => n4422, b => n4424, c => n1649, d => n3109, outb
                           => n1652);
   U2839 : aoi22 port map( a => n1652, b => mult_125_G2_ab_7_1_port, c => n4426
                           , d => n3086, outb => n4425);
   U2840 : oai22 port map( a => n4425, b => n4427, c => n1653, d => n3112, outb
                           => n1656);
   U2841 : aoi22 port map( a => n1656, b => mult_125_G2_ab_9_1_port, c => n4429
                           , d => n3089, outb => n4428);
   U2842 : oai22 port map( a => n4428, b => n4430, c => n1657, d => n3115, outb
                           => n1660);
   U2843 : aoi22 port map( a => n1660, b => mult_125_G2_ab_11_1_port, c => 
                           n4432, d => n3092, outb => n4431);
   U2844 : oai22 port map( a => n4431, b => n4433, c => n1661, d => n3118, outb
                           => n1664);
   U2845 : aoi22 port map( a => n1664, b => mult_125_G2_ab_13_1_port, c => 
                           n4435, d => n3095, outb => n4434);
   U2846 : inv port map( inb => mult_125_G2_ab_14_1_port, outb => n4436);
   U2847 : oai22 port map( a => n4434, b => n4436, c => n1665, d => n3121, outb
                           => n1668);
   U2848 : nand2 port map( a => mult_125_G2_ab_0_1_port, b => 
                           mult_125_G2_ab_1_0_port, outb => n4437);
   U2849 : aoi22 port map( a => mult_125_G2_ab_2_0_port, b => n1670, c => n4439
                           , d => n3101, outb => n4438);
   U2850 : aoi22 port map( a => n1672, b => mult_125_G2_ab_3_0_port, c => n4441
                           , d => n3102, outb => n4440);
   U2851 : inv port map( inb => mult_125_G2_ab_4_0_port, outb => n4442);
   U2852 : oai22 port map( a => n4440, b => n4442, c => n1673, d => n4443, outb
                           => n1676);
   U2853 : aoi22 port map( a => n1676, b => mult_125_G2_ab_5_0_port, c => n4445
                           , d => n3104, outb => n4444);
   U2854 : inv port map( inb => mult_125_G2_ab_6_0_port, outb => n4446);
   U2855 : oai22 port map( a => n4444, b => n4446, c => n1677, d => n4447, outb
                           => n1680);
   U2856 : aoi22 port map( a => n1680, b => mult_125_G2_ab_7_0_port, c => n4449
                           , d => n3107, outb => n4448);
   U2857 : inv port map( inb => mult_125_G2_ab_8_0_port, outb => n4450);
   U2858 : oai22 port map( a => n4448, b => n4450, c => n1681, d => n4451, outb
                           => n1684);
   U2859 : aoi22 port map( a => n1684, b => mult_125_G2_ab_9_0_port, c => n4453
                           , d => n3110, outb => n4452);
   U2860 : inv port map( inb => mult_125_G2_ab_10_0_port, outb => n4454);
   U2861 : oai22 port map( a => n4452, b => n4454, c => n1685, d => n4455, outb
                           => n1688);
   U2862 : aoi22 port map( a => n1688, b => mult_125_G2_ab_11_0_port, c => 
                           n4457, d => n3113, outb => n4456);
   U2863 : inv port map( inb => mult_125_G2_ab_12_0_port, outb => n4458);
   U2864 : oai22 port map( a => n4456, b => n4458, c => n1689, d => n4459, outb
                           => n1692);
   U2865 : aoi22 port map( a => n1692, b => mult_125_G2_ab_13_0_port, c => 
                           n4461, d => n3116, outb => n4460);
   U2866 : inv port map( inb => mult_125_G2_ab_14_0_port, outb => n4462);
   U2867 : oai22 port map( a => n4460, b => n4462, c => n1693, d => n4463, outb
                           => n1696);
   U2868 : inv port map( inb => mult_125_G2_ZB, outb => n344);
   U2869 : inv port map( inb => mult_125_G2_ZA, outb => n345);
   U2870 : nand2 port map( a => mult_125_ab_0_15_port, b => 
                           mult_125_ab_1_14_port, outb => n4464);
   U2871 : inv port map( inb => mult_125_ab_3_15_port, outb => n4465);
   U2872 : inv port map( inb => mult_125_ab_4_14_port, outb => n4466);
   U2873 : inv port map( inb => mult_125_ab_5_15_port, outb => n4467);
   U2874 : inv port map( inb => mult_125_ab_6_14_port, outb => n4468);
   U2875 : inv port map( inb => mult_125_ab_7_15_port, outb => n4469);
   U2876 : inv port map( inb => mult_125_ab_8_14_port, outb => n4470);
   U2877 : inv port map( inb => mult_125_ab_9_15_port, outb => n4471);
   U2878 : inv port map( inb => mult_125_ab_10_14_port, outb => n4472);
   U2879 : inv port map( inb => mult_125_ab_11_15_port, outb => n4473);
   U2880 : inv port map( inb => mult_125_ab_12_14_port, outb => n4474);
   U2881 : nand2 port map( a => mult_125_ab_0_14_port, b => 
                           mult_125_ab_1_13_port, outb => n1714);
   U2882 : aoi22 port map( a => mult_125_ab_2_13_port, b => n4475, c => n1712, 
                           d => n3131, outb => n1717);
   U2883 : oai22 port map( a => n1717, b => n1716, c => n4476, d => n3132, outb
                           => n1719);
   U2884 : aoi22 port map( a => n1719, b => mult_125_ab_4_13_port, c => n4478, 
                           d => n3139, outb => n4477);
   U2885 : oai22 port map( a => n4477, b => n4479, c => n1720, d => n3142, outb
                           => n1723);
   U2886 : aoi22 port map( a => n1723, b => mult_125_ab_6_13_port, c => n4481, 
                           d => n3145, outb => n4480);
   U2887 : inv port map( inb => mult_125_ab_7_13_port, outb => n4482);
   U2888 : oai22 port map( a => n4480, b => n4482, c => n1724, d => n3148, outb
                           => n1727);
   U2889 : aoi22 port map( a => n1727, b => mult_125_ab_8_13_port, c => n4484, 
                           d => n3151, outb => n4483);
   U2890 : inv port map( inb => mult_125_ab_9_13_port, outb => n4485);
   U2891 : oai22 port map( a => n4483, b => n4485, c => n1728, d => n3154, outb
                           => n1731);
   U2892 : aoi22 port map( a => n1731, b => mult_125_ab_10_13_port, c => n4487,
                           d => n3157, outb => n4486);
   U2893 : inv port map( inb => mult_125_ab_11_13_port, outb => n4488);
   U2894 : oai22 port map( a => n4486, b => n4488, c => n1732, d => n3160, outb
                           => n1735);
   U2895 : aoi22 port map( a => n1735, b => mult_125_ab_12_13_port, c => n4490,
                           d => n3163, outb => n4489);
   U2896 : inv port map( inb => mult_125_ab_13_13_port, outb => n4491);
   U2897 : oai22 port map( a => n4489, b => n4491, c => n1736, d => n3166, outb
                           => n1739);
   U2898 : aoi22 port map( a => n1739, b => mult_125_ab_14_13_port, c => n4493,
                           d => n3169, outb => n4492);
   U2899 : nand2 port map( a => mult_125_ab_0_13_port, b => 
                           mult_125_ab_1_12_port, outb => n1744);
   U2900 : aoi22 port map( a => mult_125_ab_2_12_port, b => n4495, c => n1742, 
                           d => n3134, outb => n4494);
   U2901 : oai22 port map( a => n4494, b => n4496, c => n1745, d => n3135, outb
                           => n1748);
   U2902 : aoi22 port map( a => n1748, b => mult_125_ab_4_12_port, c => n4498, 
                           d => n3177, outb => n4497);
   U2903 : aoi22 port map( a => n1750, b => mult_125_ab_5_12_port, c => n4500, 
                           d => n3137, outb => n4499);
   U2904 : inv port map( inb => mult_125_ab_6_12_port, outb => n4501);
   U2905 : oai22 port map( a => n4499, b => n4501, c => n1751, d => n3140, outb
                           => n1754);
   U2906 : aoi22 port map( a => n1754, b => mult_125_ab_7_12_port, c => n4503, 
                           d => n3143, outb => n4502);
   U2907 : inv port map( inb => mult_125_ab_8_12_port, outb => n4504);
   U2908 : oai22 port map( a => n4502, b => n4504, c => n1755, d => n3146, outb
                           => n1758);
   U2909 : aoi22 port map( a => n1758, b => mult_125_ab_9_12_port, c => n4506, 
                           d => n3149, outb => n4505);
   U2910 : inv port map( inb => mult_125_ab_10_12_port, outb => n4507);
   U2911 : oai22 port map( a => n4505, b => n4507, c => n1759, d => n3152, outb
                           => n1762);
   U2912 : aoi22 port map( a => n1762, b => mult_125_ab_11_12_port, c => n4509,
                           d => n3155, outb => n4508);
   U2913 : inv port map( inb => mult_125_ab_12_12_port, outb => n4510);
   U2914 : oai22 port map( a => n4508, b => n4510, c => n1763, d => n3158, outb
                           => n1766);
   U2915 : aoi22 port map( a => n1766, b => mult_125_ab_13_12_port, c => n4512,
                           d => n3161, outb => n4511);
   U2916 : inv port map( inb => mult_125_ab_14_12_port, outb => n4513);
   U2917 : oai22 port map( a => n4511, b => n4513, c => n1767, d => n3164, outb
                           => n1770);
   U2918 : nand2 port map( a => mult_125_ab_0_12_port, b => 
                           mult_125_ab_1_11_port, outb => n1773);
   U2919 : aoi22 port map( a => mult_125_ab_2_11_port, b => n4514, c => n1771, 
                           d => n3172, outb => n1776);
   U2920 : oai22 port map( a => n1776, b => n1775, c => n4515, d => n3173, outb
                           => n1778);
   U2921 : oai22 port map( a => n4516, b => n4517, c => n1777, d => n3183, outb
                           => n1780);
   U2922 : aoi22 port map( a => n1780, b => mult_125_ab_5_11_port, c => n4519, 
                           d => n3175, outb => n4518);
   U2923 : oai22 port map( a => n4518, b => n4520, c => n1781, d => n3186, outb
                           => n1784);
   U2924 : oai22 port map( a => n4521, b => n4522, c => n1783, d => n3189, outb
                           => n1786);
   U2925 : aoi22 port map( a => n1786, b => mult_125_ab_8_11_port, c => n4524, 
                           d => n3192, outb => n4523);
   U2926 : inv port map( inb => mult_125_ab_9_11_port, outb => n4525);
   U2927 : oai22 port map( a => n4523, b => n4525, c => n1787, d => n3195, outb
                           => n1790);
   U2928 : aoi22 port map( a => n1790, b => mult_125_ab_10_11_port, c => n4527,
                           d => n3198, outb => n4526);
   U2929 : inv port map( inb => mult_125_ab_11_11_port, outb => n4528);
   U2930 : oai22 port map( a => n4526, b => n4528, c => n1791, d => n3201, outb
                           => n1794);
   U2931 : aoi22 port map( a => n1794, b => mult_125_ab_12_11_port, c => n4530,
                           d => n3204, outb => n4529);
   U2932 : inv port map( inb => mult_125_ab_13_11_port, outb => n4531);
   U2933 : oai22 port map( a => n4529, b => n4531, c => n1795, d => n3207, outb
                           => n1798);
   U2934 : aoi22 port map( a => n1798, b => mult_125_ab_14_11_port, c => n4532,
                           d => n3210, outb => n1801);
   U2935 : nand2 port map( a => mult_125_ab_0_11_port, b => 
                           mult_125_ab_1_10_port, outb => n1804);
   U2936 : aoi22 port map( a => mult_125_ab_2_10_port, b => n4534, c => n1802, 
                           d => n3178, outb => n4533);
   U2937 : oai22 port map( a => n4533, b => n4535, c => n1805, d => n3179, outb
                           => n1808);
   U2938 : aoi22 port map( a => n1808, b => mult_125_ab_4_10_port, c => n4536, 
                           d => n3218, outb => n1811);
   U2939 : oai22 port map( a => n1811, b => n1810, c => n4537, d => n3181, outb
                           => n1813);
   U2940 : aoi22 port map( a => n1813, b => mult_125_ab_6_10_port, c => n4539, 
                           d => n3221, outb => n4538);
   U2941 : oai22 port map( a => n4538, b => n4540, c => n1814, d => n3184, outb
                           => n1817);
   U2942 : inv port map( inb => mult_125_ab_8_10_port, outb => n4541);
   U2943 : oai22 port map( a => n4542, b => n4541, c => n1816, d => n3187, outb
                           => n1819);
   U2944 : aoi22 port map( a => n1819, b => mult_125_ab_9_10_port, c => n4544, 
                           d => n3190, outb => n4543);
   U2945 : inv port map( inb => mult_125_ab_10_10_port, outb => n4545);
   U2946 : oai22 port map( a => n4543, b => n4545, c => n1820, d => n3193, outb
                           => n1823);
   U2947 : aoi22 port map( a => n1823, b => mult_125_ab_11_10_port, c => n4547,
                           d => n3196, outb => n4546);
   U2948 : inv port map( inb => mult_125_ab_12_10_port, outb => n4548);
   U2949 : oai22 port map( a => n4546, b => n4548, c => n1824, d => n3199, outb
                           => n1827);
   U2950 : aoi22 port map( a => n1827, b => mult_125_ab_13_10_port, c => n4550,
                           d => n3202, outb => n4549);
   U2951 : inv port map( inb => mult_125_ab_14_10_port, outb => n4551);
   U2952 : oai22 port map( a => n4549, b => n4551, c => n1828, d => n3205, outb
                           => n1831);
   U2953 : nand2 port map( a => mult_125_ab_0_10_port, b => 
                           mult_125_ab_1_9_port, outb => n1834);
   U2954 : aoi22 port map( a => mult_125_ab_2_9_port, b => n4553, c => n1832, d
                           => n3213, outb => n4552);
   U2955 : oai22 port map( a => n4552, b => n4554, c => n1835, d => n3214, outb
                           => n1838);
   U2956 : oai22 port map( a => n4555, b => n4556, c => n1837, d => n3227, outb
                           => n1840);
   U2957 : aoi22 port map( a => n1840, b => mult_125_ab_5_9_port, c => n4558, d
                           => n3216, outb => n4557);
   U2958 : oai22 port map( a => n4557, b => n4559, c => n1841, d => n3230, outb
                           => n1844);
   U2959 : aoi22 port map( a => n1844, b => mult_125_ab_7_9_port, c => n4561, d
                           => n3219, outb => n4560);
   U2960 : oai22 port map( a => n4560, b => n4562, c => n1845, d => n3233, outb
                           => n1848);
   U2961 : oai22 port map( a => n4563, b => n4564, c => n1847, d => n3236, outb
                           => n1850);
   U2962 : aoi22 port map( a => n1850, b => mult_125_ab_10_9_port, c => n4566, 
                           d => n3239, outb => n4565);
   U2963 : inv port map( inb => mult_125_ab_11_9_port, outb => n4567);
   U2964 : oai22 port map( a => n4565, b => n4567, c => n1851, d => n3242, outb
                           => n1854);
   U2965 : aoi22 port map( a => n1854, b => mult_125_ab_12_9_port, c => n4569, 
                           d => n3245, outb => n4568);
   U2966 : inv port map( inb => mult_125_ab_13_9_port, outb => n4570);
   U2967 : oai22 port map( a => n4568, b => n4570, c => n1855, d => n3248, outb
                           => n1858);
   U2968 : aoi22 port map( a => n1858, b => mult_125_ab_14_9_port, c => n4571, 
                           d => n3251, outb => n1861);
   U2969 : nand2 port map( a => mult_125_ab_0_9_port, b => mult_125_ab_1_8_port
                           , outb => n1864);
   U2970 : aoi22 port map( a => mult_125_ab_2_8_port, b => n4573, c => n1862, d
                           => n3222, outb => n4572);
   U2971 : oai22 port map( a => n4572, b => n4574, c => n1865, d => n3223, outb
                           => n1868);
   U2972 : oai22 port map( a => n4575, b => n4576, c => n1867, d => n3259, outb
                           => n1870);
   U2973 : oai22 port map( a => n4577, b => n4578, c => n1869, d => n3225, outb
                           => n1872);
   U2974 : aoi22 port map( a => n1872, b => mult_125_ab_6_8_port, c => n4580, d
                           => n3262, outb => n4579);
   U2975 : oai22 port map( a => n4579, b => n4581, c => n1873, d => n3228, outb
                           => n1876);
   U2976 : aoi22 port map( a => n1876, b => mult_125_ab_8_8_port, c => n4583, d
                           => n3265, outb => n4582);
   U2977 : oai22 port map( a => n4582, b => n4584, c => n1877, d => n3231, outb
                           => n1880);
   U2978 : inv port map( inb => mult_125_ab_10_8_port, outb => n4585);
   U2979 : oai22 port map( a => n4586, b => n4585, c => n1879, d => n3234, outb
                           => n1882);
   U2980 : aoi22 port map( a => n1882, b => mult_125_ab_11_8_port, c => n4588, 
                           d => n3237, outb => n4587);
   U2981 : inv port map( inb => mult_125_ab_12_8_port, outb => n4589);
   U2982 : oai22 port map( a => n4587, b => n4589, c => n1883, d => n3240, outb
                           => n1886);
   U2983 : aoi22 port map( a => n1886, b => mult_125_ab_13_8_port, c => n4591, 
                           d => n3243, outb => n4590);
   U2984 : inv port map( inb => mult_125_ab_14_8_port, outb => n4592);
   U2985 : oai22 port map( a => n4590, b => n4592, c => n1887, d => n3246, outb
                           => n1890);
   U2986 : nand2 port map( a => mult_125_ab_0_8_port, b => mult_125_ab_1_7_port
                           , outb => n1893);
   U2987 : aoi22 port map( a => mult_125_ab_2_7_port, b => n4593, c => n1891, d
                           => n3254, outb => n1896);
   U2988 : oai22 port map( a => n1896, b => n1895, c => n4594, d => n3255, outb
                           => n1898);
   U2989 : oai22 port map( a => n4595, b => n4596, c => n1897, d => n3271, outb
                           => n1900);
   U2990 : aoi22 port map( a => n1900, b => mult_125_ab_5_7_port, c => n4598, d
                           => n3257, outb => n4597);
   U2991 : oai22 port map( a => n4597, b => n4599, c => n1901, d => n3274, outb
                           => n1904);
   U2992 : aoi22 port map( a => n1904, b => mult_125_ab_7_7_port, c => n4601, d
                           => n3260, outb => n4600);
   U2993 : oai22 port map( a => n4600, b => n4602, c => n1905, d => n3277, outb
                           => n1908);
   U2994 : aoi22 port map( a => n1908, b => mult_125_ab_9_7_port, c => n4604, d
                           => n3263, outb => n4603);
   U2995 : oai22 port map( a => n4603, b => n4605, c => n1909, d => n3280, outb
                           => n1912);
   U2996 : oai22 port map( a => n4606, b => n4607, c => n1911, d => n3283, outb
                           => n1914);
   U2997 : aoi22 port map( a => n1914, b => mult_125_ab_12_7_port, c => n4609, 
                           d => n3286, outb => n4608);
   U2998 : inv port map( inb => mult_125_ab_13_7_port, outb => n4610);
   U2999 : oai22 port map( a => n4608, b => n4610, c => n1915, d => n3289, outb
                           => n1918);
   U3000 : aoi22 port map( a => n1918, b => mult_125_ab_14_7_port, c => n4611, 
                           d => n3292, outb => n1921);
   U3001 : nand2 port map( a => mult_125_ab_0_7_port, b => mult_125_ab_1_6_port
                           , outb => n1924);
   U3002 : aoi22 port map( a => mult_125_ab_2_6_port, b => n4613, c => n1922, d
                           => n3266, outb => n4612);
   U3003 : oai22 port map( a => n4612, b => n4614, c => n1925, d => n3267, outb
                           => n1928);
   U3004 : aoi22 port map( a => n1928, b => mult_125_ab_4_6_port, c => n4615, d
                           => n3300, outb => n1931);
   U3005 : oai22 port map( a => n1931, b => n1930, c => n4616, d => n3269, outb
                           => n1933);
   U3006 : aoi22 port map( a => n1933, b => mult_125_ab_6_6_port, c => n4618, d
                           => n3303, outb => n4617);
   U3007 : oai22 port map( a => n4617, b => n4619, c => n1934, d => n3272, outb
                           => n1937);
   U3008 : aoi22 port map( a => n1937, b => mult_125_ab_8_6_port, c => n4620, d
                           => n3306, outb => n1940);
   U3009 : oai22 port map( a => n1940, b => n1939, c => n4621, d => n3275, outb
                           => n1942);
   U3010 : aoi22 port map( a => n1942, b => mult_125_ab_10_6_port, c => n4623, 
                           d => n3309, outb => n4622);
   U3011 : oai22 port map( a => n4622, b => n4624, c => n1943, d => n3278, outb
                           => n1946);
   U3012 : inv port map( inb => mult_125_ab_12_6_port, outb => n4625);
   U3013 : oai22 port map( a => n4626, b => n4625, c => n1945, d => n3281, outb
                           => n1948);
   U3014 : aoi22 port map( a => n1948, b => mult_125_ab_13_6_port, c => n4628, 
                           d => n3284, outb => n4627);
   U3015 : inv port map( inb => mult_125_ab_14_6_port, outb => n4629);
   U3016 : oai22 port map( a => n4627, b => n4629, c => n1949, d => n3287, outb
                           => n1952);
   U3017 : nand2 port map( a => mult_125_ab_0_6_port, b => mult_125_ab_1_5_port
                           , outb => n1955);
   U3018 : aoi22 port map( a => mult_125_ab_2_5_port, b => n4630, c => n1953, d
                           => n3295, outb => n1958);
   U3019 : oai22 port map( a => n1958, b => n1957, c => n4631, d => n3296, outb
                           => n1960);
   U3020 : oai22 port map( a => n4632, b => n4633, c => n1959, d => n3315, outb
                           => n1962);
   U3021 : aoi22 port map( a => n1962, b => mult_125_ab_5_5_port, c => n4634, d
                           => n3298, outb => n1965);
   U3022 : oai22 port map( a => n1965, b => n1964, c => n4635, d => n3318, outb
                           => n1967);
   U3023 : aoi22 port map( a => n1967, b => mult_125_ab_7_5_port, c => n4637, d
                           => n3301, outb => n4636);
   U3024 : oai22 port map( a => n4636, b => n4638, c => n1968, d => n3321, outb
                           => n1971);
   U3025 : aoi22 port map( a => n1971, b => mult_125_ab_9_5_port, c => n4640, d
                           => n3304, outb => n4639);
   U3026 : oai22 port map( a => n4639, b => n4641, c => n1972, d => n3324, outb
                           => n1975);
   U3027 : aoi22 port map( a => n1975, b => mult_125_ab_11_5_port, c => n4643, 
                           d => n3307, outb => n4642);
   U3028 : oai22 port map( a => n4642, b => n4644, c => n1976, d => n3327, outb
                           => n1979);
   U3029 : oai22 port map( a => n4645, b => n4646, c => n1978, d => n3330, outb
                           => n1981);
   U3030 : aoi22 port map( a => n1981, b => mult_125_ab_14_5_port, c => n4647, 
                           d => n3333, outb => n1984);
   U3031 : nand2 port map( a => mult_125_ab_0_5_port, b => mult_125_ab_1_4_port
                           , outb => n1987);
   U3032 : aoi22 port map( a => mult_125_ab_2_4_port, b => n4649, c => n1985, d
                           => n3310, outb => n4648);
   U3033 : oai22 port map( a => n4648, b => n4650, c => n1988, d => n3311, outb
                           => n1991);
   U3034 : aoi22 port map( a => n1991, b => mult_125_ab_4_4_port, c => n4651, d
                           => n3341, outb => n1994);
   U3035 : oai22 port map( a => n1994, b => n1993, c => n4652, d => n3313, outb
                           => n1996);
   U3036 : aoi22 port map( a => n1996, b => mult_125_ab_6_4_port, c => n4653, d
                           => n3344, outb => n1999);
   U3037 : oai22 port map( a => n1999, b => n1998, c => n4654, d => n3316, outb
                           => n2001);
   U3038 : aoi22 port map( a => n2001, b => mult_125_ab_8_4_port, c => n4656, d
                           => n3347, outb => n4655);
   U3039 : oai22 port map( a => n4655, b => n4657, c => n2002, d => n3319, outb
                           => n2005);
   U3040 : aoi22 port map( a => n2005, b => mult_125_ab_10_4_port, c => n4658, 
                           d => n3350, outb => n2008);
   U3041 : oai22 port map( a => n2008, b => n2007, c => n4659, d => n3322, outb
                           => n2010);
   U3042 : aoi22 port map( a => n2010, b => mult_125_ab_12_4_port, c => n4661, 
                           d => n3353, outb => n4660);
   U3043 : oai22 port map( a => n4660, b => n4662, c => n2011, d => n3325, outb
                           => n2014);
   U3044 : aoi22 port map( a => n2014, b => mult_125_ab_14_4_port, c => n4663, 
                           d => n3328, outb => n2017);
   U3045 : nand2 port map( a => mult_125_ab_0_4_port, b => mult_125_ab_1_3_port
                           , outb => n2020);
   U3046 : aoi22 port map( a => mult_125_ab_2_3_port, b => n4664, c => n2018, d
                           => n3336, outb => n2023);
   U3047 : oai22 port map( a => n2023, b => n2022, c => n4665, d => n3337, outb
                           => n2025);
   U3048 : oai22 port map( a => n4666, b => n4667, c => n2024, d => n3359, outb
                           => n2027);
   U3049 : aoi22 port map( a => n2027, b => mult_125_ab_5_3_port, c => n4669, d
                           => n3339, outb => n4668);
   U3050 : oai22 port map( a => n4668, b => n4670, c => n2028, d => n3362, outb
                           => n2031);
   U3051 : aoi22 port map( a => n2031, b => mult_125_ab_7_3_port, c => n4672, d
                           => n3342, outb => n4671);
   U3052 : oai22 port map( a => n4671, b => n4673, c => n2032, d => n3365, outb
                           => n2035);
   U3053 : aoi22 port map( a => n2035, b => mult_125_ab_9_3_port, c => n4675, d
                           => n3345, outb => n4674);
   U3054 : oai22 port map( a => n4674, b => n4676, c => n2036, d => n3368, outb
                           => n2039);
   U3055 : aoi22 port map( a => n2039, b => mult_125_ab_11_3_port, c => n4678, 
                           d => n3348, outb => n4677);
   U3056 : oai22 port map( a => n4677, b => n4679, c => n2040, d => n3371, outb
                           => n2043);
   U3057 : aoi22 port map( a => n2043, b => mult_125_ab_13_3_port, c => n4681, 
                           d => n3351, outb => n4680);
   U3058 : inv port map( inb => mult_125_ab_14_3_port, outb => n4682);
   U3059 : oai22 port map( a => n4680, b => n4682, c => n2044, d => n3374, outb
                           => n2047);
   U3060 : nand2 port map( a => mult_125_ab_0_3_port, b => mult_125_ab_1_2_port
                           , outb => n2050);
   U3061 : aoi22 port map( a => mult_125_ab_2_2_port, b => n4684, c => n2048, d
                           => n3354, outb => n4683);
   U3062 : oai22 port map( a => n4683, b => n4685, c => n2051, d => n3355, outb
                           => n2054);
   U3063 : aoi22 port map( a => n2054, b => mult_125_ab_4_2_port, c => n4687, d
                           => n3382, outb => n4686);
   U3064 : oai22 port map( a => n4686, b => n4688, c => n2055, d => n3357, outb
                           => n2058);
   U3065 : aoi22 port map( a => n2058, b => mult_125_ab_6_2_port, c => n4689, d
                           => n3385, outb => n2061);
   U3066 : oai22 port map( a => n2061, b => n2060, c => n4690, d => n3360, outb
                           => n2063);
   U3067 : aoi22 port map( a => n2063, b => mult_125_ab_8_2_port, c => n4692, d
                           => n3388, outb => n4691);
   U3068 : oai22 port map( a => n4691, b => n4693, c => n2064, d => n3363, outb
                           => n2067);
   U3069 : aoi22 port map( a => n2067, b => mult_125_ab_10_2_port, c => n4695, 
                           d => n3391, outb => n4694);
   U3070 : oai22 port map( a => n4694, b => n4696, c => n2068, d => n3366, outb
                           => n2071);
   U3071 : aoi22 port map( a => n2071, b => mult_125_ab_12_2_port, c => n4698, 
                           d => n3394, outb => n4697);
   U3072 : oai22 port map( a => n4697, b => n4699, c => n2072, d => n3369, outb
                           => n2075);
   U3073 : aoi22 port map( a => n2075, b => mult_125_ab_14_2_port, c => n4701, 
                           d => n3397, outb => n4700);
   U3074 : nand2 port map( a => mult_125_ab_0_2_port, b => mult_125_ab_1_1_port
                           , outb => n2080);
   U3075 : aoi22 port map( a => mult_125_ab_2_1_port, b => n4703, c => n2078, d
                           => n3377, outb => n4702);
   U3076 : oai22 port map( a => n4702, b => n4704, c => n2081, d => n3378, outb
                           => n2084);
   U3077 : inv port map( inb => mult_125_ab_4_1_port, outb => n4705);
   U3078 : oai22 port map( a => n4706, b => n4705, c => n2083, d => n3403, outb
                           => n2086);
   U3079 : aoi22 port map( a => n2086, b => mult_125_ab_5_1_port, c => n4708, d
                           => n3380, outb => n4707);
   U3080 : oai22 port map( a => n4707, b => n4709, c => n2087, d => n3406, outb
                           => n2090);
   U3081 : aoi22 port map( a => n2090, b => mult_125_ab_7_1_port, c => n4711, d
                           => n3383, outb => n4710);
   U3082 : oai22 port map( a => n4710, b => n4712, c => n2091, d => n3409, outb
                           => n2094);
   U3083 : aoi22 port map( a => n2094, b => mult_125_ab_9_1_port, c => n4714, d
                           => n3386, outb => n4713);
   U3084 : oai22 port map( a => n4713, b => n4715, c => n2095, d => n3412, outb
                           => n2098);
   U3085 : aoi22 port map( a => n2098, b => mult_125_ab_11_1_port, c => n4717, 
                           d => n3389, outb => n4716);
   U3086 : oai22 port map( a => n4716, b => n4718, c => n2099, d => n3415, outb
                           => n2102);
   U3087 : aoi22 port map( a => n2102, b => mult_125_ab_13_1_port, c => n4720, 
                           d => n3392, outb => n4719);
   U3088 : inv port map( inb => mult_125_ab_14_1_port, outb => n4721);
   U3089 : oai22 port map( a => n4719, b => n4721, c => n2103, d => n3418, outb
                           => n2106);
   U3090 : nand2 port map( a => mult_125_ab_0_1_port, b => mult_125_ab_1_0_port
                           , outb => n4722);
   U3091 : aoi22 port map( a => mult_125_ab_2_0_port, b => n2108, c => n4724, d
                           => n3398, outb => n4723);
   U3092 : aoi22 port map( a => n2110, b => mult_125_ab_3_0_port, c => n4726, d
                           => n3399, outb => n4725);
   U3093 : inv port map( inb => mult_125_ab_4_0_port, outb => n4727);
   U3094 : oai22 port map( a => n4725, b => n4727, c => n2111, d => n4728, outb
                           => n2114);
   U3095 : aoi22 port map( a => n2114, b => mult_125_ab_5_0_port, c => n4730, d
                           => n3401, outb => n4729);
   U3096 : inv port map( inb => mult_125_ab_6_0_port, outb => n4731);
   U3097 : oai22 port map( a => n4729, b => n4731, c => n2115, d => n4732, outb
                           => n2118);
   U3098 : aoi22 port map( a => n2118, b => mult_125_ab_7_0_port, c => n4734, d
                           => n3404, outb => n4733);
   U3099 : inv port map( inb => mult_125_ab_8_0_port, outb => n4735);
   U3100 : oai22 port map( a => n4733, b => n4735, c => n2119, d => n4736, outb
                           => n2122);
   U3101 : aoi22 port map( a => n2122, b => mult_125_ab_9_0_port, c => n4738, d
                           => n3407, outb => n4737);
   U3102 : inv port map( inb => mult_125_ab_10_0_port, outb => n4739);
   U3103 : oai22 port map( a => n4737, b => n4739, c => n2123, d => n4740, outb
                           => n2126);
   U3104 : aoi22 port map( a => n2126, b => mult_125_ab_11_0_port, c => n4742, 
                           d => n3410, outb => n4741);
   U3105 : inv port map( inb => mult_125_ab_12_0_port, outb => n4743);
   U3106 : oai22 port map( a => n4741, b => n4743, c => n2127, d => n4744, outb
                           => n2130);
   U3107 : aoi22 port map( a => n2130, b => mult_125_ab_13_0_port, c => n4746, 
                           d => n3413, outb => n4745);
   U3108 : inv port map( inb => mult_125_ab_14_0_port, outb => n4747);
   U3109 : oai22 port map( a => n4745, b => n4747, c => n2131, d => n4748, outb
                           => n2134);
   U3110 : inv port map( inb => mult_125_ZB, outb => n308);
   U3111 : inv port map( inb => mult_125_ZA, outb => n309);
   U3112 : nand2 port map( a => adder_mem_array_3_0_port, b => 
                           multiplier_sigs_2_0_port, outb => n4749);
   U3113 : inv port map( inb => multiplier_sigs_2_2_port, outb => n4750);
   U3114 : inv port map( inb => adder_mem_array_3_2_port, outb => n4751);
   U3115 : inv port map( inb => multiplier_sigs_2_4_port, outb => n4752);
   U3116 : inv port map( inb => adder_mem_array_3_4_port, outb => n4753);
   U3117 : inv port map( inb => multiplier_sigs_2_6_port, outb => n4754);
   U3118 : inv port map( inb => adder_mem_array_3_6_port, outb => n4755);
   U3119 : inv port map( inb => multiplier_sigs_2_8_port, outb => n4756);
   U3120 : inv port map( inb => adder_mem_array_3_8_port, outb => n4757);
   U3121 : inv port map( inb => multiplier_sigs_2_10_port, outb => n4758);
   U3122 : inv port map( inb => adder_mem_array_3_10_port, outb => n4759);
   U3123 : inv port map( inb => multiplier_sigs_2_12_port, outb => n4760);
   U3124 : inv port map( inb => adder_mem_array_3_12_port, outb => n4761);
   U3125 : inv port map( inb => multiplier_sigs_2_14_port, outb => n4762);
   U3126 : inv port map( inb => adder_mem_array_3_14_port, outb => n4763);
   U3127 : inv port map( inb => multiplier_sigs_2_16_port, outb => n4764);
   U3128 : inv port map( inb => adder_mem_array_3_16_port, outb => n4765);
   U3129 : inv port map( inb => multiplier_sigs_2_18_port, outb => n4766);
   U3130 : inv port map( inb => adder_mem_array_3_18_port, outb => n4767);
   U3131 : inv port map( inb => multiplier_sigs_2_20_port, outb => n4768);
   U3132 : inv port map( inb => adder_mem_array_3_20_port, outb => n4769);
   U3133 : inv port map( inb => multiplier_sigs_2_22_port, outb => n4770);
   U3134 : inv port map( inb => adder_mem_array_3_22_port, outb => n4771);
   U3135 : inv port map( inb => multiplier_sigs_2_24_port, outb => n4772);
   U3136 : inv port map( inb => adder_mem_array_3_24_port, outb => n4773);
   U3137 : inv port map( inb => multiplier_sigs_2_26_port, outb => n4774);
   U3138 : inv port map( inb => adder_mem_array_3_26_port, outb => n4775);
   U3139 : nand2 port map( a => adder_mem_array_1_0_port, b => 
                           multiplier_sigs_0_0_port, outb => n4776);
   U3140 : inv port map( inb => multiplier_sigs_0_2_port, outb => n4777);
   U3141 : inv port map( inb => adder_mem_array_1_2_port, outb => n4778);
   U3142 : nand2 port map( a => adder_mem_array_2_0_port, b => 
                           multiplier_sigs_1_0_port, outb => n4779);
   U3143 : inv port map( inb => multiplier_sigs_1_2_port, outb => n4780);
   U3144 : inv port map( inb => adder_mem_array_2_2_port, outb => n4781);
   U3145 : inv port map( inb => multiplier_sigs_1_4_port, outb => n4782);
   U3146 : inv port map( inb => adder_mem_array_2_4_port, outb => n4783);
   U3147 : inv port map( inb => multiplier_sigs_1_6_port, outb => n4784);
   U3148 : inv port map( inb => adder_mem_array_2_6_port, outb => n4785);
   U3149 : inv port map( inb => multiplier_sigs_1_8_port, outb => n4786);
   U3150 : inv port map( inb => adder_mem_array_2_8_port, outb => n4787);
   U3151 : inv port map( inb => multiplier_sigs_1_10_port, outb => n4788);
   U3152 : inv port map( inb => adder_mem_array_2_10_port, outb => n4789);
   U3153 : inv port map( inb => multiplier_sigs_1_12_port, outb => n4790);
   U3154 : inv port map( inb => adder_mem_array_2_12_port, outb => n4791);
   U3155 : inv port map( inb => multiplier_sigs_1_14_port, outb => n4792);
   U3156 : inv port map( inb => adder_mem_array_2_14_port, outb => n4793);
   U3157 : inv port map( inb => multiplier_sigs_1_16_port, outb => n4794);
   U3158 : inv port map( inb => adder_mem_array_2_16_port, outb => n4795);
   U3159 : inv port map( inb => multiplier_sigs_1_18_port, outb => n4796);
   U3160 : inv port map( inb => adder_mem_array_2_18_port, outb => n4797);
   U3161 : inv port map( inb => multiplier_sigs_1_20_port, outb => n4798);
   U3162 : inv port map( inb => adder_mem_array_2_20_port, outb => n4799);
   U3163 : inv port map( inb => multiplier_sigs_1_22_port, outb => n4800);
   U3164 : inv port map( inb => adder_mem_array_2_22_port, outb => n4801);
   U3165 : inv port map( inb => multiplier_sigs_1_24_port, outb => n4802);
   U3166 : inv port map( inb => adder_mem_array_2_24_port, outb => n4803);
   U3167 : inv port map( inb => multiplier_sigs_1_26_port, outb => n4804);
   U3168 : inv port map( inb => adder_mem_array_2_26_port, outb => n4805);
   U3169 : inv port map( inb => multiplier_sigs_1_28_port, outb => n4806);
   U3170 : inv port map( inb => adder_mem_array_2_28_port, outb => n4807);
   U3171 : inv port map( inb => multiplier_sigs_1_30_port, outb => n4808);
   U3172 : inv port map( inb => adder_mem_array_2_30_port, outb => n4809);
   U3173 : inv port map( inb => multiplier_sigs_0_4_port, outb => n4810);
   U3174 : inv port map( inb => adder_mem_array_1_4_port, outb => n4811);
   U3175 : inv port map( inb => multiplier_sigs_0_6_port, outb => n4812);
   U3176 : inv port map( inb => adder_mem_array_1_6_port, outb => n4813);
   U3177 : inv port map( inb => multiplier_sigs_0_8_port, outb => n4814);
   U3178 : inv port map( inb => adder_mem_array_1_8_port, outb => n4815);
   U3179 : inv port map( inb => multiplier_sigs_0_10_port, outb => n4816);
   U3180 : inv port map( inb => adder_mem_array_1_10_port, outb => n4817);
   U3181 : inv port map( inb => multiplier_sigs_0_12_port, outb => n4818);
   U3182 : inv port map( inb => adder_mem_array_1_12_port, outb => n4819);
   U3183 : inv port map( inb => multiplier_sigs_0_14_port, outb => n4820);
   U3184 : inv port map( inb => adder_mem_array_1_14_port, outb => n4821);
   U3185 : inv port map( inb => multiplier_sigs_0_16_port, outb => n4822);
   U3186 : inv port map( inb => adder_mem_array_1_16_port, outb => n4823);
   U3187 : inv port map( inb => multiplier_sigs_0_18_port, outb => n4824);
   U3188 : inv port map( inb => adder_mem_array_1_18_port, outb => n4825);
   U3189 : inv port map( inb => multiplier_sigs_0_20_port, outb => n4826);
   U3190 : inv port map( inb => adder_mem_array_1_20_port, outb => n4827);
   U3191 : inv port map( inb => multiplier_sigs_0_22_port, outb => n4828);
   U3192 : inv port map( inb => adder_mem_array_1_22_port, outb => n4829);
   U3193 : inv port map( inb => multiplier_sigs_0_24_port, outb => n4830);
   U3194 : inv port map( inb => adder_mem_array_1_24_port, outb => n4831);
   U3195 : inv port map( inb => multiplier_sigs_0_26_port, outb => n4832);
   U3196 : inv port map( inb => adder_mem_array_1_26_port, outb => n4833);
   U3197 : inv port map( inb => multiplier_sigs_0_28_port, outb => n4834);
   U3198 : inv port map( inb => adder_mem_array_1_28_port, outb => n4835);
   U3199 : inv port map( inb => multiplier_sigs_0_30_port, outb => n4836);
   U3200 : inv port map( inb => adder_mem_array_1_30_port, outb => n4837);
   U3201 : inv port map( inb => multiplier_sigs_2_28_port, outb => n4838);
   U3202 : inv port map( inb => adder_mem_array_3_28_port, outb => n4839);
   U3203 : inv port map( inb => multiplier_sigs_2_30_port, outb => n4840);
   U3204 : inv port map( inb => adder_mem_array_3_30_port, outb => n4841);
   U3205 : xor2 port map( a => mult_125_G4_ab_0_1_port, b => 
                           mult_125_G4_ab_1_0_port, outb => 
                           multiplier_sigs_3_1_port);
   U3206 : xor2 port map( a => n3885, b => n4842, outb => mult_125_G4_A1_8_port
                           );
   U3207 : xor2 port map( a => n3881, b => n4843, outb => mult_125_G4_A1_6_port
                           );
   U3208 : xor2 port map( a => n3877, b => n4844, outb => mult_125_G4_A1_4_port
                           );
   U3209 : xor2 port map( a => n3873, b => n4845, outb => mult_125_G4_A1_2_port
                           );
   U3210 : xor2 port map( a => n243, b => n244, outb => mult_125_G4_A1_27_port)
                           ;
   U3211 : xor2 port map( a => n247, b => n248, outb => mult_125_G4_A1_25_port)
                           ;
   U3212 : xor2 port map( a => n251, b => n252, outb => mult_125_G4_A1_23_port)
                           ;
   U3213 : xor2 port map( a => n255, b => n256, outb => mult_125_G4_A1_21_port)
                           ;
   U3214 : xor2 port map( a => n259, b => n260, outb => mult_125_G4_A1_19_port)
                           ;
   U3215 : xor2 port map( a => n263, b => n264, outb => mult_125_G4_A1_17_port)
                           ;
   U3216 : xor2 port map( a => n268, b => n269, outb => mult_125_G4_A1_15_port)
                           ;
   U3217 : xor2 port map( a => n270, b => n271, outb => mult_125_G4_A1_14_port)
                           ;
   U3218 : xor2 port map( a => n3893, b => n4846, outb => 
                           mult_125_G4_A1_12_port);
   U3219 : xor2 port map( a => n3889, b => n4847, outb => 
                           mult_125_G4_A1_10_port);
   U3220 : xor2 port map( a => n2507, b => n4848, outb => mult_125_G4_A1_0_port
                           );
   U3221 : xor2 port map( a => n4170, b => n4849, outb => mult_125_G3_A1_8_port
                           );
   U3222 : xor2 port map( a => n4166, b => n4850, outb => mult_125_G3_A1_6_port
                           );
   U3223 : xor2 port map( a => n4162, b => n4851, outb => mult_125_G3_A1_4_port
                           );
   U3224 : xor2 port map( a => n4158, b => n4852, outb => mult_125_G3_A1_2_port
                           );
   U3225 : xor2 port map( a => n351, b => n352, outb => mult_125_G3_A1_27_port)
                           ;
   U3226 : xor2 port map( a => n355, b => n356, outb => mult_125_G3_A1_25_port)
                           ;
   U3227 : xor2 port map( a => n359, b => n360, outb => mult_125_G3_A1_23_port)
                           ;
   U3228 : xor2 port map( a => n363, b => n364, outb => mult_125_G3_A1_21_port)
                           ;
   U3229 : xor2 port map( a => n367, b => n368, outb => mult_125_G3_A1_19_port)
                           ;
   U3230 : xor2 port map( a => n371, b => n372, outb => mult_125_G3_A1_17_port)
                           ;
   U3231 : xor2 port map( a => n376, b => n377, outb => mult_125_G3_A1_15_port)
                           ;
   U3232 : xor2 port map( a => n378, b => n379, outb => mult_125_G3_A1_14_port)
                           ;
   U3233 : xor2 port map( a => n4178, b => n4853, outb => 
                           mult_125_G3_A1_12_port);
   U3234 : xor2 port map( a => n4174, b => n4854, outb => 
                           mult_125_G3_A1_10_port);
   U3235 : xor2 port map( a => n2804, b => n4855, outb => mult_125_G3_A1_0_port
                           );
   U3236 : xor2 port map( a => n4455, b => n4856, outb => mult_125_G2_A1_8_port
                           );
   U3237 : xor2 port map( a => n4451, b => n4857, outb => mult_125_G2_A1_6_port
                           );
   U3238 : xor2 port map( a => n4447, b => n4858, outb => mult_125_G2_A1_4_port
                           );
   U3239 : xor2 port map( a => n4443, b => n4859, outb => mult_125_G2_A1_2_port
                           );
   U3240 : xor2 port map( a => n315, b => n316, outb => mult_125_G2_A1_27_port)
                           ;
   U3241 : xor2 port map( a => n319, b => n320, outb => mult_125_G2_A1_25_port)
                           ;
   U3242 : xor2 port map( a => n323, b => n324, outb => mult_125_G2_A1_23_port)
                           ;
   U3243 : xor2 port map( a => n327, b => n328, outb => mult_125_G2_A1_21_port)
                           ;
   U3244 : xor2 port map( a => n331, b => n332, outb => mult_125_G2_A1_19_port)
                           ;
   U3245 : xor2 port map( a => n335, b => n336, outb => mult_125_G2_A1_17_port)
                           ;
   U3246 : xor2 port map( a => n340, b => n341, outb => mult_125_G2_A1_15_port)
                           ;
   U3247 : xor2 port map( a => n342, b => n343, outb => mult_125_G2_A1_14_port)
                           ;
   U3248 : xor2 port map( a => n4463, b => n4860, outb => 
                           mult_125_G2_A1_12_port);
   U3249 : xor2 port map( a => n4459, b => n4861, outb => 
                           mult_125_G2_A1_10_port);
   U3250 : xor2 port map( a => n3101, b => n4862, outb => mult_125_G2_A1_0_port
                           );
   U3251 : xor2 port map( a => n4740, b => n4863, outb => mult_125_A1_8_port);
   U3252 : xor2 port map( a => n4736, b => n4864, outb => mult_125_A1_6_port);
   U3253 : xor2 port map( a => n4732, b => n4865, outb => mult_125_A1_4_port);
   U3254 : xor2 port map( a => n4728, b => n4866, outb => mult_125_A1_2_port);
   U3255 : xor2 port map( a => n279, b => n280, outb => mult_125_A1_27_port);
   U3256 : xor2 port map( a => n283, b => n284, outb => mult_125_A1_25_port);
   U3257 : xor2 port map( a => n287, b => n288, outb => mult_125_A1_23_port);
   U3258 : xor2 port map( a => n291, b => n292, outb => mult_125_A1_21_port);
   U3259 : xor2 port map( a => n295, b => n296, outb => mult_125_A1_19_port);
   U3260 : xor2 port map( a => n299, b => n300, outb => mult_125_A1_17_port);
   U3261 : xor2 port map( a => n304, b => n305, outb => mult_125_A1_15_port);
   U3262 : xor2 port map( a => n306, b => n307, outb => mult_125_A1_14_port);
   U3263 : xor2 port map( a => n4748, b => n4867, outb => mult_125_A1_12_port);
   U3264 : xor2 port map( a => n4744, b => n4868, outb => mult_125_A1_10_port);
   U3265 : xor2 port map( a => n3398, b => n4869, outb => mult_125_A1_0_port);
   U3266 : xor2 port map( a => n3426, b => n4870, outb => N73);
   U3267 : xor2 port map( a => adder_mem_array_3_0_port, b => 
                           multiplier_sigs_2_0_port, outb => N72);
   U3268 : xor2 port map( a => n3447, b => n4871, outb => N7);
   U3269 : xor2 port map( a => adder_mem_array_1_0_port, b => 
                           multiplier_sigs_0_0_port, outb => N6);
   U3270 : xor2 port map( a => n3484, b => n4872, outb => N40);
   U3271 : xor2 port map( a => adder_mem_array_2_0_port, b => 
                           multiplier_sigs_1_0_port, outb => N39);
   U3272 : xor2 port map( a => mult_125_G4_QA, b => mult_125_G4_QB, outb => 
                           n2239);
   U3273 : xor2 port map( a => mult_125_G4_ab_3_14_port, b => 
                           mult_125_G4_ab_2_15_port, outb => n4873);
   U3274 : xor2 port map( a => mult_125_G4_ab_5_14_port, b => 
                           mult_125_G4_ab_4_15_port, outb => n4874);
   U3275 : xor2 port map( a => mult_125_G4_ab_7_14_port, b => 
                           mult_125_G4_ab_6_15_port, outb => n4875);
   U3276 : xor2 port map( a => mult_125_G4_ab_9_14_port, b => 
                           mult_125_G4_ab_8_15_port, outb => n4876);
   U3277 : xor2 port map( a => mult_125_G4_ab_11_14_port, b => 
                           mult_125_G4_ab_10_15_port, outb => n4877);
   U3278 : xor2 port map( a => mult_125_G4_ab_13_14_port, b => 
                           mult_125_G4_ab_12_15_port, outb => n4878);
   U3279 : xor2 port map( a => mult_125_G4_ab_15_14_port, b => 
                           mult_125_G4_ab_14_15_port, outb => n4879);
   U3280 : xor2 port map( a => mult_125_G4_ab_10_0_port, b => n3882, outb => 
                           n4842);
   U3281 : xor2 port map( a => mult_125_G4_ab_8_0_port, b => n3878, outb => 
                           n4843);
   U3282 : xor2 port map( a => mult_125_G4_ab_6_0_port, b => n3874, outb => 
                           n4844);
   U3283 : xor2 port map( a => n3872, b => n798, outb => n4845);
   U3284 : xor2 port map( a => mult_125_G4_ab_14_0_port, b => n3890, outb => 
                           n4846);
   U3285 : xor2 port map( a => mult_125_G4_ab_12_0_port, b => n3886, outb => 
                           n4847);
   U3286 : xor2 port map( a => n794, b => mult_125_G4_ab_2_0_port, outb => 
                           n4848);
   U3287 : xor2 port map( a => mult_125_G3_QA, b => mult_125_G3_QB, outb => 
                           n2536);
   U3288 : xor2 port map( a => mult_125_G3_ab_3_14_port, b => 
                           mult_125_G3_ab_2_15_port, outb => n4880);
   U3289 : xor2 port map( a => mult_125_G3_ab_5_14_port, b => 
                           mult_125_G3_ab_4_15_port, outb => n4881);
   U3290 : xor2 port map( a => mult_125_G3_ab_7_14_port, b => 
                           mult_125_G3_ab_6_15_port, outb => n4882);
   U3291 : xor2 port map( a => mult_125_G3_ab_9_14_port, b => 
                           mult_125_G3_ab_8_15_port, outb => n4883);
   U3292 : xor2 port map( a => mult_125_G3_ab_11_14_port, b => 
                           mult_125_G3_ab_10_15_port, outb => n4884);
   U3293 : xor2 port map( a => mult_125_G3_ab_13_14_port, b => 
                           mult_125_G3_ab_12_15_port, outb => n4885);
   U3294 : xor2 port map( a => mult_125_G3_ab_15_14_port, b => 
                           mult_125_G3_ab_14_15_port, outb => n4886);
   U3295 : xor2 port map( a => mult_125_G3_ab_10_0_port, b => n4167, outb => 
                           n4849);
   U3296 : xor2 port map( a => mult_125_G3_ab_8_0_port, b => n4163, outb => 
                           n4850);
   U3297 : xor2 port map( a => mult_125_G3_ab_6_0_port, b => n4159, outb => 
                           n4851);
   U3298 : xor2 port map( a => n4157, b => n1236, outb => n4852);
   U3299 : xor2 port map( a => mult_125_G3_ab_14_0_port, b => n4175, outb => 
                           n4853);
   U3300 : xor2 port map( a => mult_125_G3_ab_12_0_port, b => n4171, outb => 
                           n4854);
   U3301 : xor2 port map( a => n1232, b => mult_125_G3_ab_2_0_port, outb => 
                           n4855);
   U3302 : xor2 port map( a => mult_125_G2_QA, b => mult_125_G2_QB, outb => 
                           n2833);
   U3303 : xor2 port map( a => mult_125_G2_ab_3_14_port, b => 
                           mult_125_G2_ab_2_15_port, outb => n4887);
   U3304 : xor2 port map( a => mult_125_G2_ab_5_14_port, b => 
                           mult_125_G2_ab_4_15_port, outb => n4888);
   U3305 : xor2 port map( a => mult_125_G2_ab_7_14_port, b => 
                           mult_125_G2_ab_6_15_port, outb => n4889);
   U3306 : xor2 port map( a => mult_125_G2_ab_9_14_port, b => 
                           mult_125_G2_ab_8_15_port, outb => n4890);
   U3307 : xor2 port map( a => mult_125_G2_ab_11_14_port, b => 
                           mult_125_G2_ab_10_15_port, outb => n4891);
   U3308 : xor2 port map( a => mult_125_G2_ab_13_14_port, b => 
                           mult_125_G2_ab_12_15_port, outb => n4892);
   U3309 : xor2 port map( a => mult_125_G2_ab_15_14_port, b => 
                           mult_125_G2_ab_14_15_port, outb => n4893);
   U3310 : xor2 port map( a => mult_125_G2_ab_10_0_port, b => n4452, outb => 
                           n4856);
   U3311 : xor2 port map( a => mult_125_G2_ab_8_0_port, b => n4448, outb => 
                           n4857);
   U3312 : xor2 port map( a => mult_125_G2_ab_6_0_port, b => n4444, outb => 
                           n4858);
   U3313 : xor2 port map( a => n4442, b => n1674, outb => n4859);
   U3314 : xor2 port map( a => mult_125_G2_ab_14_0_port, b => n4460, outb => 
                           n4860);
   U3315 : xor2 port map( a => mult_125_G2_ab_12_0_port, b => n4456, outb => 
                           n4861);
   U3316 : xor2 port map( a => n1670, b => mult_125_G2_ab_2_0_port, outb => 
                           n4862);
   U3317 : xor2 port map( a => mult_125_QA, b => mult_125_QB, outb => n3130);
   U3318 : xor2 port map( a => mult_125_ab_3_14_port, b => 
                           mult_125_ab_2_15_port, outb => n4894);
   U3319 : xor2 port map( a => mult_125_ab_5_14_port, b => 
                           mult_125_ab_4_15_port, outb => n4895);
   U3320 : xor2 port map( a => mult_125_ab_7_14_port, b => 
                           mult_125_ab_6_15_port, outb => n4896);
   U3321 : xor2 port map( a => mult_125_ab_9_14_port, b => 
                           mult_125_ab_8_15_port, outb => n4897);
   U3322 : xor2 port map( a => mult_125_ab_11_14_port, b => 
                           mult_125_ab_10_15_port, outb => n4898);
   U3323 : xor2 port map( a => mult_125_ab_13_14_port, b => 
                           mult_125_ab_12_15_port, outb => n4899);
   U3324 : xor2 port map( a => mult_125_ab_15_14_port, b => 
                           mult_125_ab_14_15_port, outb => n4900);
   U3325 : xor2 port map( a => mult_125_ab_10_0_port, b => n4737, outb => n4863
                           );
   U3326 : xor2 port map( a => mult_125_ab_8_0_port, b => n4733, outb => n4864)
                           ;
   U3327 : xor2 port map( a => mult_125_ab_6_0_port, b => n4729, outb => n4865)
                           ;
   U3328 : xor2 port map( a => n4727, b => n2112, outb => n4866);
   U3329 : xor2 port map( a => mult_125_ab_14_0_port, b => n4745, outb => n4867
                           );
   U3330 : xor2 port map( a => mult_125_ab_12_0_port, b => n4741, outb => n4868
                           );
   U3331 : xor2 port map( a => n2108, b => mult_125_ab_2_0_port, outb => n4869)
                           ;
   U3332 : xor2 port map( a => adder_mem_array_3_27_port, b => 
                           multiplier_sigs_2_27_port, outb => n3428);
   U3333 : xor2 port map( a => adder_mem_array_3_25_port, b => 
                           multiplier_sigs_2_25_port, outb => n3432);
   U3334 : xor2 port map( a => adder_mem_array_3_23_port, b => 
                           multiplier_sigs_2_23_port, outb => n3436);
   U3335 : xor2 port map( a => adder_mem_array_3_21_port, b => 
                           multiplier_sigs_2_21_port, outb => n3440);
   U3336 : xor2 port map( a => adder_mem_array_3_19_port, b => 
                           multiplier_sigs_2_19_port, outb => n3444);
   U3337 : xor2 port map( a => adder_mem_array_1_3_port, b => 
                           multiplier_sigs_0_3_port, outb => n3449);
   U3338 : xor2 port map( a => adder_mem_array_3_17_port, b => 
                           multiplier_sigs_2_17_port, outb => n3451);
   U3339 : xor2 port map( a => adder_mem_array_3_15_port, b => 
                           multiplier_sigs_2_15_port, outb => n3455);
   U3340 : xor2 port map( a => adder_mem_array_3_13_port, b => 
                           multiplier_sigs_2_13_port, outb => n3459);
   U3341 : xor2 port map( a => adder_mem_array_3_11_port, b => 
                           multiplier_sigs_2_11_port, outb => n3463);
   U3342 : xor2 port map( a => adder_mem_array_3_9_port, b => 
                           multiplier_sigs_2_9_port, outb => n3467);
   U3343 : xor2 port map( a => adder_mem_array_3_7_port, b => 
                           multiplier_sigs_2_7_port, outb => n3473);
   U3344 : xor2 port map( a => adder_mem_array_3_5_port, b => 
                           multiplier_sigs_2_5_port, outb => n3477);
   U3345 : xor2 port map( a => adder_mem_array_3_3_port, b => 
                           multiplier_sigs_2_3_port, outb => n3481);
   U3346 : xor2 port map( a => n2137, b => adder_mem_array_3_1_port, outb => 
                           n4870);
   U3347 : xor2 port map( a => adder_mem_array_2_31_port, b => 
                           multiplier_sigs_1_31_port, outb => n3486);
   U3348 : xor2 port map( a => n2164, b => adder_mem_array_1_1_port, outb => 
                           n4871);
   U3349 : xor2 port map( a => adder_mem_array_2_29_port, b => 
                           multiplier_sigs_1_29_port, outb => n3490);
   U3350 : xor2 port map( a => adder_mem_array_2_27_port, b => 
                           multiplier_sigs_1_27_port, outb => n3494);
   U3351 : xor2 port map( a => adder_mem_array_2_25_port, b => 
                           multiplier_sigs_1_25_port, outb => n3498);
   U3352 : xor2 port map( a => adder_mem_array_2_23_port, b => 
                           multiplier_sigs_1_23_port, outb => n3502);
   U3353 : xor2 port map( a => adder_mem_array_2_21_port, b => 
                           multiplier_sigs_1_21_port, outb => n3506);
   U3354 : xor2 port map( a => adder_mem_array_2_19_port, b => 
                           multiplier_sigs_1_19_port, outb => n3510);
   U3355 : xor2 port map( a => adder_mem_array_2_17_port, b => 
                           multiplier_sigs_1_17_port, outb => n3514);
   U3356 : xor2 port map( a => adder_mem_array_2_15_port, b => 
                           multiplier_sigs_1_15_port, outb => n3518);
   U3357 : xor2 port map( a => adder_mem_array_2_13_port, b => 
                           multiplier_sigs_1_13_port, outb => n3522);
   U3358 : xor2 port map( a => adder_mem_array_2_11_port, b => 
                           multiplier_sigs_1_11_port, outb => n3526);
   U3359 : xor2 port map( a => adder_mem_array_2_9_port, b => 
                           multiplier_sigs_1_9_port, outb => n3530);
   U3360 : xor2 port map( a => adder_mem_array_2_7_port, b => 
                           multiplier_sigs_1_7_port, outb => n3534);
   U3361 : xor2 port map( a => adder_mem_array_2_5_port, b => 
                           multiplier_sigs_1_5_port, outb => n3538);
   U3362 : xor2 port map( a => adder_mem_array_2_3_port, b => 
                           multiplier_sigs_1_3_port, outb => n3542);
   U3363 : xor2 port map( a => n2167, b => adder_mem_array_2_1_port, outb => 
                           n4872);
   U3364 : xor2 port map( a => adder_mem_array_1_31_port, b => 
                           multiplier_sigs_0_31_port, outb => n3546);
   U3365 : xor2 port map( a => adder_mem_array_1_29_port, b => 
                           multiplier_sigs_0_29_port, outb => n3550);
   U3366 : xor2 port map( a => adder_mem_array_1_27_port, b => 
                           multiplier_sigs_0_27_port, outb => n3554);
   U3367 : xor2 port map( a => adder_mem_array_1_25_port, b => 
                           multiplier_sigs_0_25_port, outb => n3558);
   U3368 : xor2 port map( a => adder_mem_array_1_23_port, b => 
                           multiplier_sigs_0_23_port, outb => n3562);
   U3369 : xor2 port map( a => adder_mem_array_1_21_port, b => 
                           multiplier_sigs_0_21_port, outb => n3566);
   U3370 : xor2 port map( a => adder_mem_array_1_19_port, b => 
                           multiplier_sigs_0_19_port, outb => n3570);
   U3371 : xor2 port map( a => adder_mem_array_1_17_port, b => 
                           multiplier_sigs_0_17_port, outb => n3574);
   U3372 : xor2 port map( a => adder_mem_array_1_15_port, b => 
                           multiplier_sigs_0_15_port, outb => n3578);
   U3373 : xor2 port map( a => adder_mem_array_1_13_port, b => 
                           multiplier_sigs_0_13_port, outb => n3582);
   U3374 : xor2 port map( a => adder_mem_array_1_11_port, b => 
                           multiplier_sigs_0_11_port, outb => n3586);
   U3375 : xor2 port map( a => adder_mem_array_1_9_port, b => 
                           multiplier_sigs_0_9_port, outb => n3590);
   U3376 : xor2 port map( a => adder_mem_array_1_7_port, b => 
                           multiplier_sigs_0_7_port, outb => n3594);
   U3377 : xor2 port map( a => adder_mem_array_1_5_port, b => 
                           multiplier_sigs_0_5_port, outb => n3598);
   U3378 : xor2 port map( a => adder_mem_array_3_31_port, b => 
                           multiplier_sigs_2_31_port, outb => n3600);
   U3379 : xor2 port map( a => adder_mem_array_3_29_port, b => 
                           multiplier_sigs_2_29_port, outb => n3604);
   U3380 : oai22 port map( a => n4902, b => n4903, c => n384, d => n3609, outb 
                           => n4901);
   U3381 : aoi22 port map( a => mult_125_G4_ab_2_15_port, b => 
                           mult_125_G4_ab_3_14_port, c => n4901, d => n4905, 
                           outb => n4904);
   U3382 : oai22 port map( a => n3610, b => n3611, c => n4904, d => n386, outb 
                           => n4906);
   U3383 : aoi22 port map( a => mult_125_G4_ab_4_15_port, b => 
                           mult_125_G4_ab_5_14_port, c => n4906, d => n4908, 
                           outb => n4907);
   U3384 : oai22 port map( a => n3612, b => n3613, c => n4907, d => n388, outb 
                           => n4909);
   U3385 : aoi22 port map( a => mult_125_G4_ab_6_15_port, b => 
                           mult_125_G4_ab_7_14_port, c => n4909, d => n4911, 
                           outb => n4910);
   U3386 : oai22 port map( a => n3614, b => n3615, c => n4910, d => n390, outb 
                           => n4912);
   U3387 : aoi22 port map( a => mult_125_G4_ab_8_15_port, b => 
                           mult_125_G4_ab_9_14_port, c => n4912, d => n4914, 
                           outb => n4913);
   U3388 : oai22 port map( a => n3616, b => n3617, c => n4913, d => n392, outb 
                           => n4915);
   U3389 : aoi22 port map( a => mult_125_G4_ab_10_15_port, b => 
                           mult_125_G4_ab_11_14_port, c => n4915, d => n4917, 
                           outb => n4916);
   U3390 : oai22 port map( a => n3618, b => n3619, c => n4916, d => n394, outb 
                           => n4918);
   U3391 : aoi22 port map( a => mult_125_G4_ab_12_15_port, b => 
                           mult_125_G4_ab_13_14_port, c => n4918, d => n4920, 
                           outb => n4919);
   U3392 : aoi22 port map( a => mult_125_G4_ab_13_15_port, b => 
                           mult_125_G4_ab_14_14_port, c => n4922, d => n4923, 
                           outb => n4921);
   U3393 : aoi22 port map( a => mult_125_G4_ab_14_15_port, b => 
                           mult_125_G4_ab_15_14_port, c => n4924, d => n4925, 
                           outb => n241);
   U3394 : inv port map( inb => n3637, outb => n427);
   U3395 : aoi22 port map( a => n427, b => mult_125_G4_ab_15_13_port, c => 
                           n4926, d => n2280, outb => n243);
   U3396 : aoi22 port map( a => n456, b => mult_125_G4_ab_15_12_port, c => 
                           n4927, d => n2276, outb => n245);
   U3397 : oai22 port map( a => n487, b => n486, c => n4929, d => n2321, outb 
                           => n4928);
   U3398 : inv port map( inb => n503, outb => n3687);
   U3399 : aoi22 port map( a => n517, b => mult_125_G4_ab_15_10_port, c => 
                           n4930, d => n2317, outb => n249);
   U3400 : oai22 port map( a => n547, b => n546, c => n4932, d => n2362, outb 
                           => n4931);
   U3401 : inv port map( inb => n566, outb => n3731);
   U3402 : aoi22 port map( a => n576, b => mult_125_G4_ab_15_8_port, c => n4933
                           , d => n2358, outb => n253);
   U3403 : oai22 port map( a => n607, b => n606, c => n4935, d => n2403, outb 
                           => n4934);
   U3404 : inv port map( inb => n632, outb => n3771);
   U3405 : aoi22 port map( a => n638, b => mult_125_G4_ab_15_6_port, c => n4936
                           , d => n2399, outb => n257);
   U3406 : oai22 port map( a => n670, b => n669, c => n4938, d => n2444, outb 
                           => n4937);
   U3407 : aoi22 port map( a => n4939, b => mult_125_G4_ab_15_4_port, c => n701
                           , d => n2440, outb => n261);
   U3408 : aoi22 port map( a => n733, b => mult_125_G4_ab_15_3_port, c => n4940
                           , d => n2485, outb => n263);
   U3409 : oai22 port map( a => n3845, b => n4941, c => n762, d => n2481, outb 
                           => n266);
   U3410 : aoi22 port map( a => n792, b => mult_125_G4_ab_15_1_port, c => n4942
                           , d => n2504, outb => n268);
   U3411 : aoi22 port map( a => n820, b => mult_125_G4_ab_15_0_port, c => n4943
                           , d => n4944, outb => n270);
   U3412 : xor2 port map( a => n4901, b => n4873, outb => n2248);
   U3413 : xor2 port map( a => n4945, b => n4904, outb => n2251);
   U3414 : xor2 port map( a => n4906, b => n4874, outb => n2254);
   U3415 : xor2 port map( a => n4946, b => n4907, outb => n2257);
   U3416 : xor2 port map( a => n4909, b => n4875, outb => n2260);
   U3417 : xor2 port map( a => n4947, b => n4910, outb => n2263);
   U3418 : xor2 port map( a => n4912, b => n4876, outb => n2266);
   U3419 : xor2 port map( a => n4948, b => n4913, outb => n2269);
   U3420 : xor2 port map( a => n4915, b => n4877, outb => n2272);
   U3421 : xor2 port map( a => n4949, b => n4916, outb => n2275);
   U3422 : xor2 port map( a => n4918, b => n4878, outb => n2278);
   U3423 : xor2 port map( a => n4950, b => n4922, outb => n2280);
   U3424 : xor2 port map( a => n4921, b => n4879, outb => n244);
   U3425 : xor2 port map( a => n4951, b => n2241, outb => n2286);
   U3426 : xor2 port map( a => n4952, b => n2244, outb => n2292);
   U3427 : xor2 port map( a => n4953, b => n2246, outb => n2295);
   U3428 : xor2 port map( a => n4954, b => n2249, outb => n2298);
   U3429 : xor2 port map( a => n4955, b => n2252, outb => n2301);
   U3430 : xor2 port map( a => n4956, b => n2255, outb => n2304);
   U3431 : xor2 port map( a => n4957, b => n2258, outb => n2307);
   U3432 : xor2 port map( a => n4958, b => n2261, outb => n2310);
   U3433 : xor2 port map( a => n4959, b => n2264, outb => n2313);
   U3434 : xor2 port map( a => n4960, b => n2267, outb => n2316);
   U3435 : xor2 port map( a => n4961, b => n2270, outb => n2319);
   U3436 : xor2 port map( a => n4962, b => n2273, outb => n2321);
   U3437 : xor2 port map( a => n4963, b => n2276, outb => n248);
   U3438 : xor2 port map( a => n4964, b => n2282, outb => n2327);
   U3439 : xor2 port map( a => n4965, b => n2284, outb => n2330);
   U3440 : xor2 port map( a => n4966, b => n2288, outb => n2336);
   U3441 : xor2 port map( a => n4967, b => n2290, outb => n2339);
   U3442 : xor2 port map( a => n4968, b => n2293, outb => n2342);
   U3443 : xor2 port map( a => n4969, b => n2296, outb => n2345);
   U3444 : xor2 port map( a => n4970, b => n2299, outb => n2348);
   U3445 : xor2 port map( a => n4971, b => n2302, outb => n2351);
   U3446 : xor2 port map( a => n4972, b => n2305, outb => n2354);
   U3447 : xor2 port map( a => n4973, b => n2308, outb => n2357);
   U3448 : xor2 port map( a => n4974, b => n2311, outb => n2360);
   U3449 : xor2 port map( a => n4975, b => n2314, outb => n2362);
   U3450 : xor2 port map( a => n4976, b => n2317, outb => n252);
   U3451 : xor2 port map( a => n4977, b => n2323, outb => n2368);
   U3452 : xor2 port map( a => n4978, b => n2325, outb => n2371);
   U3453 : xor2 port map( a => n4979, b => n2328, outb => n2374);
   U3454 : xor2 port map( a => n4980, b => n2332, outb => n2380);
   U3455 : xor2 port map( a => n4981, b => n2334, outb => n2383);
   U3456 : xor2 port map( a => n4982, b => n2337, outb => n2386);
   U3457 : xor2 port map( a => n4983, b => n2340, outb => n2389);
   U3458 : xor2 port map( a => n4984, b => n2343, outb => n2392);
   U3459 : xor2 port map( a => n4985, b => n2346, outb => n2395);
   U3460 : xor2 port map( a => n4986, b => n2349, outb => n2398);
   U3461 : xor2 port map( a => n4987, b => n2352, outb => n2401);
   U3462 : xor2 port map( a => n4988, b => n2355, outb => n2403);
   U3463 : xor2 port map( a => n4989, b => n2358, outb => n256);
   U3464 : xor2 port map( a => n4990, b => n2364, outb => n2409);
   U3465 : xor2 port map( a => n4991, b => n2366, outb => n2412);
   U3466 : xor2 port map( a => n4992, b => n2369, outb => n2415);
   U3467 : xor2 port map( a => n4993, b => n2372, outb => n2418);
   U3468 : xor2 port map( a => n4994, b => n2376, outb => n2424);
   U3469 : xor2 port map( a => n4995, b => n2378, outb => n2427);
   U3470 : xor2 port map( a => n4996, b => n2381, outb => n2430);
   U3471 : xor2 port map( a => n4997, b => n2384, outb => n2433);
   U3472 : xor2 port map( a => n4998, b => n2387, outb => n2436);
   U3473 : xor2 port map( a => n4999, b => n2390, outb => n2439);
   U3474 : xor2 port map( a => n5000, b => n2393, outb => n2442);
   U3475 : xor2 port map( a => n5001, b => n2396, outb => n2444);
   U3476 : xor2 port map( a => n5002, b => n2399, outb => n260);
   U3477 : xor2 port map( a => n5003, b => n2405, outb => n2450);
   U3478 : xor2 port map( a => n5004, b => n2407, outb => n2453);
   U3479 : xor2 port map( a => n5005, b => n2410, outb => n2456);
   U3480 : xor2 port map( a => n5006, b => n2413, outb => n2459);
   U3481 : xor2 port map( a => n5007, b => n2416, outb => n2462);
   U3482 : xor2 port map( a => n5008, b => n2420, outb => n2468);
   U3483 : xor2 port map( a => n5009, b => n2422, outb => n2471);
   U3484 : xor2 port map( a => n5010, b => n2425, outb => n2474);
   U3485 : xor2 port map( a => n5011, b => n2428, outb => n2477);
   U3486 : xor2 port map( a => n5012, b => n2431, outb => n2480);
   U3487 : xor2 port map( a => n5013, b => n2434, outb => n2483);
   U3488 : xor2 port map( a => n5014, b => n2437, outb => n2485);
   U3489 : xor2 port map( a => n5015, b => n2440, outb => n264);
   U3490 : xor2 port map( a => n5016, b => n2446, outb => n2491);
   U3491 : xor2 port map( a => n5017, b => n2448, outb => n2494);
   U3492 : xor2 port map( a => n5018, b => n2451, outb => n2497);
   U3493 : xor2 port map( a => n5019, b => n2454, outb => n2500);
   U3494 : xor2 port map( a => n5020, b => n2457, outb => n2503);
   U3495 : xor2 port map( a => n5021, b => n2460, outb => n2506);
   U3496 : xor2 port map( a => n5022, b => n2464, outb => n2512);
   U3497 : xor2 port map( a => n5023, b => n2466, outb => n2515);
   U3498 : xor2 port map( a => n5024, b => n2469, outb => n2518);
   U3499 : xor2 port map( a => n5025, b => n2472, outb => n2521);
   U3500 : xor2 port map( a => n5026, b => n2475, outb => n2524);
   U3501 : xor2 port map( a => n5027, b => n2478, outb => n2527);
   U3502 : xor2 port map( a => n5028, b => n2481, outb => n269);
   U3503 : xor2 port map( a => n5029, b => n2487, outb => n3873);
   U3504 : xor2 port map( a => n5030, b => n2489, outb => n3877);
   U3505 : xor2 port map( a => n5031, b => n2492, outb => n3881);
   U3506 : xor2 port map( a => n5032, b => n2495, outb => n3885);
   U3507 : xor2 port map( a => n5033, b => n2498, outb => n3889);
   U3508 : xor2 port map( a => n5034, b => n2501, outb => n3893);
   U3509 : inv port map( inb => n2525, outb => n4944);
   U3510 : xor2 port map( a => n5035, b => n2504, outb => n271);
   U3511 : xor2 port map( a => n5036, b => n2525, outb => n275);
   U3512 : xor2 port map( a => n3609, b => mult_125_G4_ab_2_14_port, outb => 
                           n2242);
   U3513 : xor2 port map( a => n3610, b => n3611, outb => n4945);
   U3514 : xor2 port map( a => n3612, b => n3613, outb => n4946);
   U3515 : xor2 port map( a => n3614, b => n3615, outb => n4947);
   U3516 : xor2 port map( a => n3616, b => n3617, outb => n4948);
   U3517 : xor2 port map( a => n3618, b => n3619, outb => n4949);
   U3518 : xor2 port map( a => mult_125_G4_ab_13_15_port, b => 
                           mult_125_G4_ab_14_14_port, outb => n4950);
   U3519 : xor2 port map( a => n3620, b => n399, outb => n2245);
   U3520 : xor2 port map( a => mult_125_G4_ab_3_13_port, b => n403, outb => 
                           n4951);
   U3521 : xor2 port map( a => mult_125_G4_ab_4_13_port, b => n405, outb => 
                           n2247);
   U3522 : xor2 port map( a => mult_125_G4_ab_5_13_port, b => n407, outb => 
                           n2250);
   U3523 : xor2 port map( a => mult_125_G4_ab_6_13_port, b => n409, outb => 
                           n2253);
   U3524 : xor2 port map( a => n3627, b => n3625, outb => n2256);
   U3525 : xor2 port map( a => mult_125_G4_ab_8_13_port, b => n413, outb => 
                           n2259);
   U3526 : xor2 port map( a => n3630, b => n3628, outb => n2262);
   U3527 : xor2 port map( a => mult_125_G4_ab_10_13_port, b => n417, outb => 
                           n2265);
   U3528 : xor2 port map( a => n3633, b => n3631, outb => n2268);
   U3529 : xor2 port map( a => mult_125_G4_ab_12_13_port, b => n421, outb => 
                           n2271);
   U3530 : xor2 port map( a => n3636, b => n3634, outb => n2274);
   U3531 : xor2 port map( a => mult_125_G4_ab_14_13_port, b => n425, outb => 
                           n2277);
   U3532 : xor2 port map( a => mult_125_G4_ab_15_13_port, b => n3637, outb => 
                           n2279);
   U3533 : xor2 port map( a => n430, b => mult_125_G4_ab_2_12_port, outb => 
                           n2283);
   U3534 : xor2 port map( a => n3641, b => n3639, outb => n4952);
   U3535 : xor2 port map( a => mult_125_G4_ab_4_12_port, b => n434, outb => 
                           n2285);
   U3536 : xor2 port map( a => mult_125_G4_ab_5_12_port, b => n3642, outb => 
                           n4953);
   U3537 : xor2 port map( a => n3646, b => n3644, outb => n4954);
   U3538 : xor2 port map( a => mult_125_G4_ab_7_12_port, b => n440, outb => 
                           n4955);
   U3539 : xor2 port map( a => n3649, b => n3647, outb => n4956);
   U3540 : xor2 port map( a => mult_125_G4_ab_9_12_port, b => n444, outb => 
                           n4957);
   U3541 : xor2 port map( a => n3652, b => n3650, outb => n4958);
   U3542 : xor2 port map( a => mult_125_G4_ab_11_12_port, b => n448, outb => 
                           n4959);
   U3543 : xor2 port map( a => n3655, b => n3653, outb => n4960);
   U3544 : xor2 port map( a => mult_125_G4_ab_13_12_port, b => n452, outb => 
                           n4961);
   U3545 : xor2 port map( a => n3658, b => n3656, outb => n4962);
   U3546 : xor2 port map( a => n5037, b => n456, outb => n4963);
   U3547 : xor2 port map( a => n459, b => mult_125_G4_ab_2_11_port, outb => 
                           n2289);
   U3548 : xor2 port map( a => mult_125_G4_ab_3_11_port, b => n462, outb => 
                           n4964);
   U3549 : xor2 port map( a => n3662, b => n3661, outb => n2291);
   U3550 : xor2 port map( a => mult_125_G4_ab_5_11_port, b => n466, outb => 
                           n4965);
   U3551 : xor2 port map( a => mult_125_G4_ab_6_11_port, b => n468, outb => 
                           n2294);
   U3552 : xor2 port map( a => n3667, b => n3666, outb => n2297);
   U3553 : xor2 port map( a => mult_125_G4_ab_8_11_port, b => n472, outb => 
                           n2300);
   U3554 : xor2 port map( a => n3670, b => n3668, outb => n2303);
   U3555 : xor2 port map( a => mult_125_G4_ab_10_11_port, b => n476, outb => 
                           n2306);
   U3556 : xor2 port map( a => n3673, b => n3671, outb => n2309);
   U3557 : xor2 port map( a => mult_125_G4_ab_12_11_port, b => n480, outb => 
                           n2312);
   U3558 : xor2 port map( a => n3676, b => n3674, outb => n2315);
   U3559 : xor2 port map( a => mult_125_G4_ab_14_11_port, b => n484, outb => 
                           n2318);
   U3560 : xor2 port map( a => n486, b => n487, outb => n2320);
   U3561 : xor2 port map( a => n490, b => mult_125_G4_ab_2_10_port, outb => 
                           n2324);
   U3562 : xor2 port map( a => n3680, b => n3678, outb => n4966);
   U3563 : xor2 port map( a => mult_125_G4_ab_4_10_port, b => n494, outb => 
                           n2326);
   U3564 : xor2 port map( a => n496, b => n497, outb => n4967);
   U3565 : xor2 port map( a => mult_125_G4_ab_6_10_port, b => n499, outb => 
                           n2329);
   U3566 : xor2 port map( a => mult_125_G4_ab_7_10_port, b => n501, outb => 
                           n4968);
   U3567 : xor2 port map( a => n3686, b => n3687, outb => n4969);
   U3568 : xor2 port map( a => mult_125_G4_ab_9_10_port, b => n505, outb => 
                           n4970);
   U3569 : xor2 port map( a => n3690, b => n3688, outb => n4971);
   U3570 : xor2 port map( a => mult_125_G4_ab_11_10_port, b => n509, outb => 
                           n4972);
   U3571 : xor2 port map( a => n3693, b => n3691, outb => n4973);
   U3572 : xor2 port map( a => mult_125_G4_ab_13_10_port, b => n513, outb => 
                           n4974);
   U3573 : xor2 port map( a => n3696, b => n3694, outb => n4975);
   U3574 : xor2 port map( a => n5038, b => n517, outb => n4976);
   U3575 : xor2 port map( a => n520, b => mult_125_G4_ab_2_9_port, outb => 
                           n2333);
   U3576 : xor2 port map( a => n3699, b => n3697, outb => n4977);
   U3577 : xor2 port map( a => mult_125_G4_ab_4_9_port, b => n524, outb => 
                           n2335);
   U3578 : xor2 port map( a => mult_125_G4_ab_5_9_port, b => n526, outb => 
                           n4978);
   U3579 : xor2 port map( a => mult_125_G4_ab_6_9_port, b => n528, outb => 
                           n2338);
   U3580 : xor2 port map( a => mult_125_G4_ab_7_9_port, b => n530, outb => 
                           n4979);
   U3581 : xor2 port map( a => n3707, b => n3705, outb => n2341);
   U3582 : xor2 port map( a => n3709, b => n3708, outb => n2344);
   U3583 : xor2 port map( a => mult_125_G4_ab_10_9_port, b => n536, outb => 
                           n2347);
   U3584 : xor2 port map( a => n3712, b => n3710, outb => n2350);
   U3585 : xor2 port map( a => mult_125_G4_ab_12_9_port, b => n540, outb => 
                           n2353);
   U3586 : xor2 port map( a => n3715, b => n3713, outb => n2356);
   U3587 : xor2 port map( a => mult_125_G4_ab_14_9_port, b => n544, outb => 
                           n2359);
   U3588 : xor2 port map( a => n546, b => n547, outb => n2361);
   U3589 : xor2 port map( a => n550, b => mult_125_G4_ab_2_8_port, outb => 
                           n2365);
   U3590 : xor2 port map( a => n3719, b => n3717, outb => n4980);
   U3591 : xor2 port map( a => n3721, b => n554, outb => n2367);
   U3592 : xor2 port map( a => n3723, b => n3722, outb => n4981);
   U3593 : xor2 port map( a => mult_125_G4_ab_6_8_port, b => n558, outb => 
                           n2370);
   U3594 : xor2 port map( a => n3726, b => n3724, outb => n4982);
   U3595 : xor2 port map( a => mult_125_G4_ab_8_8_port, b => n562, outb => 
                           n2373);
   U3596 : xor2 port map( a => mult_125_G4_ab_9_8_port, b => n564, outb => 
                           n4983);
   U3597 : xor2 port map( a => n3730, b => n3731, outb => n4984);
   U3598 : xor2 port map( a => mult_125_G4_ab_11_8_port, b => n568, outb => 
                           n4985);
   U3599 : xor2 port map( a => n3734, b => n3732, outb => n4986);
   U3600 : xor2 port map( a => mult_125_G4_ab_13_8_port, b => n572, outb => 
                           n4987);
   U3601 : xor2 port map( a => n3737, b => n3735, outb => n4988);
   U3602 : xor2 port map( a => n5039, b => n576, outb => n4989);
   U3603 : xor2 port map( a => n579, b => mult_125_G4_ab_2_7_port, outb => 
                           n2377);
   U3604 : xor2 port map( a => mult_125_G4_ab_3_7_port, b => n582, outb => 
                           n4990);
   U3605 : xor2 port map( a => n3741, b => n3740, outb => n2379);
   U3606 : xor2 port map( a => mult_125_G4_ab_5_7_port, b => n586, outb => 
                           n4991);
   U3607 : xor2 port map( a => n3744, b => n3742, outb => n2382);
   U3608 : xor2 port map( a => mult_125_G4_ab_7_7_port, b => n590, outb => 
                           n4992);
   U3609 : xor2 port map( a => n3747, b => n3745, outb => n2385);
   U3610 : xor2 port map( a => mult_125_G4_ab_9_7_port, b => n594, outb => 
                           n4993);
   U3611 : xor2 port map( a => n3750, b => n3748, outb => n2388);
   U3612 : xor2 port map( a => n3752, b => n3751, outb => n2391);
   U3613 : xor2 port map( a => mult_125_G4_ab_12_7_port, b => n600, outb => 
                           n2394);
   U3614 : xor2 port map( a => n3755, b => n3753, outb => n2397);
   U3615 : xor2 port map( a => mult_125_G4_ab_14_7_port, b => n604, outb => 
                           n2400);
   U3616 : xor2 port map( a => n606, b => n607, outb => n2402);
   U3617 : xor2 port map( a => n610, b => mult_125_G4_ab_2_6_port, outb => 
                           n2406);
   U3618 : xor2 port map( a => n3759, b => n3757, outb => n4994);
   U3619 : xor2 port map( a => mult_125_G4_ab_4_6_port, b => n614, outb => 
                           n2408);
   U3620 : xor2 port map( a => n616, b => n617, outb => n4995);
   U3621 : xor2 port map( a => mult_125_G4_ab_6_6_port, b => n619, outb => 
                           n2411);
   U3622 : xor2 port map( a => n3764, b => n3762, outb => n4996);
   U3623 : xor2 port map( a => mult_125_G4_ab_8_6_port, b => n623, outb => 
                           n2414);
   U3624 : xor2 port map( a => n625, b => n626, outb => n4997);
   U3625 : xor2 port map( a => mult_125_G4_ab_10_6_port, b => n628, outb => 
                           n2417);
   U3626 : xor2 port map( a => mult_125_G4_ab_11_6_port, b => n630, outb => 
                           n4998);
   U3627 : xor2 port map( a => n3770, b => n3771, outb => n4999);
   U3628 : xor2 port map( a => mult_125_G4_ab_13_6_port, b => n634, outb => 
                           n5000);
   U3629 : xor2 port map( a => n3774, b => n3772, outb => n5001);
   U3630 : xor2 port map( a => n5040, b => n638, outb => n5002);
   U3631 : xor2 port map( a => n641, b => mult_125_G4_ab_2_5_port, outb => 
                           n2421);
   U3632 : xor2 port map( a => mult_125_G4_ab_3_5_port, b => n644, outb => 
                           n5003);
   U3633 : xor2 port map( a => mult_125_G4_ab_4_5_port, b => n646, outb => 
                           n2423);
   U3634 : xor2 port map( a => mult_125_G4_ab_5_5_port, b => n648, outb => 
                           n5004);
   U3635 : xor2 port map( a => n650, b => n651, outb => n2426);
   U3636 : xor2 port map( a => mult_125_G4_ab_7_5_port, b => n653, outb => 
                           n5005);
   U3637 : xor2 port map( a => mult_125_G4_ab_8_5_port, b => n655, outb => 
                           n2429);
   U3638 : xor2 port map( a => mult_125_G4_ab_9_5_port, b => n657, outb => 
                           n5006);
   U3639 : xor2 port map( a => n3786, b => n3784, outb => n2432);
   U3640 : xor2 port map( a => mult_125_G4_ab_11_5_port, b => n661, outb => 
                           n5007);
   U3641 : xor2 port map( a => n3789, b => n3787, outb => n2435);
   U3642 : xor2 port map( a => n3791, b => n665, outb => n2438);
   U3643 : xor2 port map( a => mult_125_G4_ab_14_5_port, b => n667, outb => 
                           n2441);
   U3644 : xor2 port map( a => n669, b => n670, outb => n2443);
   U3645 : xor2 port map( a => n673, b => mult_125_G4_ab_2_4_port, outb => 
                           n2447);
   U3646 : xor2 port map( a => n3795, b => n3793, outb => n5008);
   U3647 : xor2 port map( a => mult_125_G4_ab_4_4_port, b => n677, outb => 
                           n2449);
   U3648 : xor2 port map( a => n679, b => n680, outb => n5009);
   U3649 : xor2 port map( a => mult_125_G4_ab_6_4_port, b => n682, outb => 
                           n2452);
   U3650 : xor2 port map( a => n684, b => n685, outb => n5010);
   U3651 : xor2 port map( a => mult_125_G4_ab_8_4_port, b => n687, outb => 
                           n2455);
   U3652 : xor2 port map( a => mult_125_G4_ab_9_4_port, b => n689, outb => 
                           n5011);
   U3653 : xor2 port map( a => mult_125_G4_ab_10_4_port, b => n691, outb => 
                           n2458);
   U3654 : xor2 port map( a => n693, b => n694, outb => n5012);
   U3655 : xor2 port map( a => mult_125_G4_ab_12_4_port, b => n696, outb => 
                           n2461);
   U3656 : xor2 port map( a => mult_125_G4_ab_13_4_port, b => n698, outb => 
                           n5013);
   U3657 : xor2 port map( a => mult_125_G4_ab_14_4_port, b => n700, outb => 
                           n5014);
   U3658 : xor2 port map( a => mult_125_G4_ab_15_4_port, b => n703, outb => 
                           n5015);
   U3659 : xor2 port map( a => n706, b => mult_125_G4_ab_2_3_port, outb => 
                           n2465);
   U3660 : xor2 port map( a => mult_125_G4_ab_3_3_port, b => n709, outb => 
                           n5016);
   U3661 : xor2 port map( a => mult_125_G4_ab_4_3_port, b => n711, outb => 
                           n2467);
   U3662 : xor2 port map( a => mult_125_G4_ab_5_3_port, b => n713, outb => 
                           n5017);
   U3663 : xor2 port map( a => mult_125_G4_ab_6_3_port, b => n715, outb => 
                           n2470);
   U3664 : xor2 port map( a => mult_125_G4_ab_7_3_port, b => n717, outb => 
                           n5018);
   U3665 : xor2 port map( a => mult_125_G4_ab_8_3_port, b => n719, outb => 
                           n2473);
   U3666 : xor2 port map( a => mult_125_G4_ab_9_3_port, b => n721, outb => 
                           n5019);
   U3667 : xor2 port map( a => mult_125_G4_ab_10_3_port, b => n723, outb => 
                           n2476);
   U3668 : xor2 port map( a => mult_125_G4_ab_11_3_port, b => n725, outb => 
                           n5020);
   U3669 : xor2 port map( a => n3824, b => n3822, outb => n2479);
   U3670 : xor2 port map( a => mult_125_G4_ab_13_3_port, b => n729, outb => 
                           n5021);
   U3671 : xor2 port map( a => mult_125_G4_ab_14_3_port, b => n731, outb => 
                           n2482);
   U3672 : xor2 port map( a => mult_125_G4_ab_15_3_port, b => n733, outb => 
                           n2484);
   U3673 : xor2 port map( a => n736, b => mult_125_G4_ab_2_2_port, outb => 
                           n2488);
   U3674 : xor2 port map( a => n3830, b => n3828, outb => n5022);
   U3675 : xor2 port map( a => mult_125_G4_ab_4_2_port, b => n740, outb => 
                           n2490);
   U3676 : xor2 port map( a => mult_125_G4_ab_5_2_port, b => n742, outb => 
                           n5023);
   U3677 : xor2 port map( a => mult_125_G4_ab_6_2_port, b => n744, outb => 
                           n2493);
   U3678 : xor2 port map( a => n746, b => n747, outb => n5024);
   U3679 : xor2 port map( a => mult_125_G4_ab_8_2_port, b => n749, outb => 
                           n2496);
   U3680 : xor2 port map( a => mult_125_G4_ab_9_2_port, b => n751, outb => 
                           n5025);
   U3681 : xor2 port map( a => mult_125_G4_ab_10_2_port, b => n753, outb => 
                           n2499);
   U3682 : xor2 port map( a => mult_125_G4_ab_11_2_port, b => n755, outb => 
                           n5026);
   U3683 : xor2 port map( a => mult_125_G4_ab_12_2_port, b => n757, outb => 
                           n2502);
   U3684 : xor2 port map( a => mult_125_G4_ab_13_2_port, b => n759, outb => 
                           n5027);
   U3685 : xor2 port map( a => mult_125_G4_ab_14_2_port, b => n761, outb => 
                           n2505);
   U3686 : xor2 port map( a => n4941, b => n3845, outb => n5028);
   U3687 : xor2 port map( a => n3848, b => mult_125_G4_ab_2_1_port, outb => 
                           n2509);
   U3688 : xor2 port map( a => n3849, b => n3847, outb => n5029);
   U3689 : xor2 port map( a => mult_125_G4_ab_4_1_port, b => n3851, outb => 
                           n2511);
   U3690 : xor2 port map( a => mult_125_G4_ab_5_1_port, b => n772, outb => 
                           n5041);
   U3691 : xor2 port map( a => n3854, b => n774, outb => n2514);
   U3692 : xor2 port map( a => n5042, b => n776, outb => n5031);
   U3693 : xor2 port map( a => mult_125_G4_ab_8_1_port, b => n3855, outb => 
                           n2517);
   U3694 : xor2 port map( a => n5043, b => n780, outb => n5032);
   U3695 : xor2 port map( a => n3860, b => n782, outb => n2520);
   U3696 : xor2 port map( a => n5044, b => n784, outb => n5033);
   U3697 : xor2 port map( a => n3863, b => n786, outb => n2523);
   U3698 : xor2 port map( a => n5045, b => n788, outb => n5034);
   U3699 : xor2 port map( a => n3866, b => n3864, outb => n2526);
   U3700 : xor2 port map( a => n5046, b => n792, outb => n5035);
   U3701 : xor2 port map( a => mult_125_G4_ab_15_0_port, b => n820, outb => 
                           n5036);
   U3702 : xor2 port map( a => mult_125_G4_ab_11_0_port, b => n812, outb => 
                           n2528);
   U3703 : xor2 port map( a => mult_125_G4_ab_9_0_port, b => n808, outb => 
                           n2529);
   U3704 : xor2 port map( a => mult_125_G4_ab_7_0_port, b => n804, outb => 
                           n2530);
   U3705 : xor2 port map( a => mult_125_G4_ab_5_0_port, b => n800, outb => 
                           n2531);
   U3706 : xor2 port map( a => mult_125_G4_ab_3_0_port, b => n796, outb => 
                           n2532);
   U3707 : xor2 port map( a => n272, b => mult_125_G4_ZA, outb => n2533);
   U3708 : xor2 port map( a => mult_125_G4_ab_13_0_port, b => n816, outb => 
                           n2534);
   U3709 : oai22 port map( a => n5048, b => n5049, c => n822, d => n3894, outb 
                           => n5047);
   U3710 : aoi22 port map( a => mult_125_G3_ab_2_15_port, b => 
                           mult_125_G3_ab_3_14_port, c => n5047, d => n5051, 
                           outb => n5050);
   U3711 : oai22 port map( a => n3895, b => n3896, c => n5050, d => n824, outb 
                           => n5052);
   U3712 : aoi22 port map( a => mult_125_G3_ab_4_15_port, b => 
                           mult_125_G3_ab_5_14_port, c => n5052, d => n5054, 
                           outb => n5053);
   U3713 : oai22 port map( a => n3897, b => n3898, c => n5053, d => n826, outb 
                           => n5055);
   U3714 : aoi22 port map( a => mult_125_G3_ab_6_15_port, b => 
                           mult_125_G3_ab_7_14_port, c => n5055, d => n5057, 
                           outb => n5056);
   U3715 : oai22 port map( a => n3899, b => n3900, c => n5056, d => n828, outb 
                           => n5058);
   U3716 : aoi22 port map( a => mult_125_G3_ab_8_15_port, b => 
                           mult_125_G3_ab_9_14_port, c => n5058, d => n5060, 
                           outb => n5059);
   U3717 : oai22 port map( a => n3901, b => n3902, c => n5059, d => n830, outb 
                           => n5061);
   U3718 : aoi22 port map( a => mult_125_G3_ab_10_15_port, b => 
                           mult_125_G3_ab_11_14_port, c => n5061, d => n5063, 
                           outb => n5062);
   U3719 : oai22 port map( a => n3903, b => n3904, c => n5062, d => n832, outb 
                           => n5064);
   U3720 : aoi22 port map( a => mult_125_G3_ab_12_15_port, b => 
                           mult_125_G3_ab_13_14_port, c => n5064, d => n5066, 
                           outb => n5065);
   U3721 : aoi22 port map( a => mult_125_G3_ab_13_15_port, b => 
                           mult_125_G3_ab_14_14_port, c => n5068, d => n5069, 
                           outb => n5067);
   U3722 : aoi22 port map( a => mult_125_G3_ab_14_15_port, b => 
                           mult_125_G3_ab_15_14_port, c => n5070, d => n5071, 
                           outb => n349);
   U3723 : inv port map( inb => n3922, outb => n865);
   U3724 : aoi22 port map( a => n865, b => mult_125_G3_ab_15_13_port, c => 
                           n5072, d => n2577, outb => n351);
   U3725 : aoi22 port map( a => n894, b => mult_125_G3_ab_15_12_port, c => 
                           n5073, d => n2573, outb => n353);
   U3726 : oai22 port map( a => n925, b => n924, c => n5075, d => n2618, outb 
                           => n5074);
   U3727 : inv port map( inb => n941, outb => n3972);
   U3728 : aoi22 port map( a => n955, b => mult_125_G3_ab_15_10_port, c => 
                           n5076, d => n2614, outb => n357);
   U3729 : oai22 port map( a => n985, b => n984, c => n5078, d => n2659, outb 
                           => n5077);
   U3730 : inv port map( inb => n1004, outb => n4016);
   U3731 : aoi22 port map( a => n1014, b => mult_125_G3_ab_15_8_port, c => 
                           n5079, d => n2655, outb => n361);
   U3732 : oai22 port map( a => n1045, b => n1044, c => n5081, d => n2700, outb
                           => n5080);
   U3733 : inv port map( inb => n1070, outb => n4056);
   U3734 : aoi22 port map( a => n1076, b => mult_125_G3_ab_15_6_port, c => 
                           n5082, d => n2696, outb => n365);
   U3735 : oai22 port map( a => n1108, b => n1107, c => n5084, d => n2741, outb
                           => n5083);
   U3736 : aoi22 port map( a => n5085, b => mult_125_G3_ab_15_4_port, c => 
                           n1139, d => n2737, outb => n369);
   U3737 : aoi22 port map( a => n1171, b => mult_125_G3_ab_15_3_port, c => 
                           n5086, d => n2782, outb => n371);
   U3738 : oai22 port map( a => n4130, b => n5087, c => n1200, d => n2778, outb
                           => n374);
   U3739 : aoi22 port map( a => n1230, b => mult_125_G3_ab_15_1_port, c => 
                           n5088, d => n2801, outb => n376);
   U3740 : aoi22 port map( a => n1258, b => mult_125_G3_ab_15_0_port, c => 
                           n5089, d => n5090, outb => n378);
   U3741 : aoi22 port map( a => adder_mem_array_3_1_port, b => n2137, c => 
                           n5091, d => n3426, outb => n3483);
   U3742 : oai22 port map( a => n4750, b => n4751, c => n3483, d => n2138, outb
                           => n3480);
   U3743 : aoi22 port map( a => multiplier_sigs_2_3_port, b => 
                           adder_mem_array_3_3_port, c => n3480, d => n5092, 
                           outb => n3479);
   U3744 : oai22 port map( a => n4752, b => n4753, c => n3479, d => n2140, outb
                           => n3476);
   U3745 : aoi22 port map( a => multiplier_sigs_2_5_port, b => 
                           adder_mem_array_3_5_port, c => n3476, d => n5093, 
                           outb => n3475);
   U3746 : oai22 port map( a => n4754, b => n4755, c => n3475, d => n2142, outb
                           => n3472);
   U3747 : aoi22 port map( a => multiplier_sigs_2_7_port, b => 
                           adder_mem_array_3_7_port, c => n3472, d => n5094, 
                           outb => n3469);
   U3748 : oai22 port map( a => n4756, b => n4757, c => n3469, d => n2144, outb
                           => n3466);
   U3749 : aoi22 port map( a => multiplier_sigs_2_9_port, b => 
                           adder_mem_array_3_9_port, c => n3466, d => n5095, 
                           outb => n3465);
   U3750 : oai22 port map( a => n4758, b => n4759, c => n3465, d => n2146, outb
                           => n3462);
   U3751 : aoi22 port map( a => multiplier_sigs_2_11_port, b => 
                           adder_mem_array_3_11_port, c => n3462, d => n5096, 
                           outb => n3461);
   U3752 : oai22 port map( a => n4760, b => n4761, c => n3461, d => n2148, outb
                           => n3458);
   U3753 : aoi22 port map( a => multiplier_sigs_2_13_port, b => 
                           adder_mem_array_3_13_port, c => n3458, d => n5097, 
                           outb => n3457);
   U3754 : oai22 port map( a => n4762, b => n4763, c => n3457, d => n2150, outb
                           => n3454);
   U3755 : aoi22 port map( a => multiplier_sigs_2_15_port, b => 
                           adder_mem_array_3_15_port, c => n3454, d => n5098, 
                           outb => n3453);
   U3756 : oai22 port map( a => n4764, b => n4765, c => n3453, d => n2152, outb
                           => n3450);
   U3757 : aoi22 port map( a => multiplier_sigs_2_17_port, b => 
                           adder_mem_array_3_17_port, c => n3450, d => n5099, 
                           outb => n3446);
   U3758 : oai22 port map( a => n4766, b => n4767, c => n3446, d => n2154, outb
                           => n3443);
   U3759 : aoi22 port map( a => multiplier_sigs_2_19_port, b => 
                           adder_mem_array_3_19_port, c => n3443, d => n5100, 
                           outb => n3442);
   U3760 : oai22 port map( a => n4768, b => n4769, c => n3442, d => n2156, outb
                           => n3439);
   U3761 : aoi22 port map( a => multiplier_sigs_2_21_port, b => 
                           adder_mem_array_3_21_port, c => n3439, d => n5101, 
                           outb => n3438);
   U3762 : oai22 port map( a => n4770, b => n4771, c => n3438, d => n2158, outb
                           => n3435);
   U3763 : aoi22 port map( a => multiplier_sigs_2_23_port, b => 
                           adder_mem_array_3_23_port, c => n3435, d => n5102, 
                           outb => n3434);
   U3764 : oai22 port map( a => n4772, b => n4773, c => n3434, d => n2160, outb
                           => n3431);
   U3765 : aoi22 port map( a => multiplier_sigs_2_25_port, b => 
                           adder_mem_array_3_25_port, c => n3431, d => n5103, 
                           outb => n3430);
   U3766 : oai22 port map( a => n4774, b => n4775, c => n3430, d => n2162, outb
                           => n3427);
   U3767 : aoi22 port map( a => adder_mem_array_3_27_port, b => 
                           multiplier_sigs_2_27_port, c => n3427, d => n5104, 
                           outb => n3606);
   U3768 : oai22 port map( a => n4838, b => n4839, c => n3606, d => n2232, outb
                           => n3603);
   U3769 : aoi22 port map( a => multiplier_sigs_2_29_port, b => 
                           adder_mem_array_3_29_port, c => n3603, d => n5105, 
                           outb => n3602);
   U3770 : oai22 port map( a => n4840, b => n4841, c => n3602, d => n2234, outb
                           => n2237);
   U3771 : nand2 port map( a => n5106, b => n5107, outb => n2236);
   U3772 : xor2 port map( a => n5047, b => n4880, outb => n2545);
   U3773 : xor2 port map( a => n5108, b => n5050, outb => n2548);
   U3774 : xor2 port map( a => n5052, b => n4881, outb => n2551);
   U3775 : xor2 port map( a => n5109, b => n5053, outb => n2554);
   U3776 : xor2 port map( a => n5055, b => n4882, outb => n2557);
   U3777 : xor2 port map( a => n5110, b => n5056, outb => n2560);
   U3778 : xor2 port map( a => n5058, b => n4883, outb => n2563);
   U3779 : xor2 port map( a => n5111, b => n5059, outb => n2566);
   U3780 : xor2 port map( a => n5061, b => n4884, outb => n2569);
   U3781 : xor2 port map( a => n5112, b => n5062, outb => n2572);
   U3782 : xor2 port map( a => n5064, b => n4885, outb => n2575);
   U3783 : xor2 port map( a => n5113, b => n5068, outb => n2577);
   U3784 : xor2 port map( a => n5067, b => n4886, outb => n352);
   U3785 : xor2 port map( a => n5114, b => n2538, outb => n2583);
   U3786 : xor2 port map( a => n5115, b => n2541, outb => n2589);
   U3787 : xor2 port map( a => n5116, b => n2543, outb => n2592);
   U3788 : xor2 port map( a => n5117, b => n2546, outb => n2595);
   U3789 : xor2 port map( a => n5118, b => n2549, outb => n2598);
   U3790 : xor2 port map( a => n5119, b => n2552, outb => n2601);
   U3791 : xor2 port map( a => n5120, b => n2555, outb => n2604);
   U3792 : xor2 port map( a => n5121, b => n2558, outb => n2607);
   U3793 : xor2 port map( a => n5122, b => n2561, outb => n2610);
   U3794 : xor2 port map( a => n5123, b => n2564, outb => n2613);
   U3795 : xor2 port map( a => n5124, b => n2567, outb => n2616);
   U3796 : xor2 port map( a => n5125, b => n2570, outb => n2618);
   U3797 : xor2 port map( a => n5126, b => n2573, outb => n356);
   U3798 : xor2 port map( a => n5127, b => n2579, outb => n2624);
   U3799 : xor2 port map( a => n5128, b => n2581, outb => n2627);
   U3800 : xor2 port map( a => n5129, b => n2585, outb => n2633);
   U3801 : xor2 port map( a => n5130, b => n2587, outb => n2636);
   U3802 : xor2 port map( a => n5131, b => n2590, outb => n2639);
   U3803 : xor2 port map( a => n5132, b => n2593, outb => n2642);
   U3804 : xor2 port map( a => n5133, b => n2596, outb => n2645);
   U3805 : xor2 port map( a => n5134, b => n2599, outb => n2648);
   U3806 : xor2 port map( a => n5135, b => n2602, outb => n2651);
   U3807 : xor2 port map( a => n5136, b => n2605, outb => n2654);
   U3808 : xor2 port map( a => n5137, b => n2608, outb => n2657);
   U3809 : xor2 port map( a => n5138, b => n2611, outb => n2659);
   U3810 : xor2 port map( a => n5139, b => n2614, outb => n360);
   U3811 : xor2 port map( a => n5140, b => n2620, outb => n2665);
   U3812 : xor2 port map( a => n5141, b => n2622, outb => n2668);
   U3813 : xor2 port map( a => n5142, b => n2625, outb => n2671);
   U3814 : xor2 port map( a => n5143, b => n2629, outb => n2677);
   U3815 : xor2 port map( a => n5144, b => n2631, outb => n2680);
   U3816 : xor2 port map( a => n5145, b => n2634, outb => n2683);
   U3817 : xor2 port map( a => n5146, b => n2637, outb => n2686);
   U3818 : xor2 port map( a => n5147, b => n2640, outb => n2689);
   U3819 : xor2 port map( a => n5148, b => n2643, outb => n2692);
   U3820 : xor2 port map( a => n5149, b => n2646, outb => n2695);
   U3821 : xor2 port map( a => n5150, b => n2649, outb => n2698);
   U3822 : xor2 port map( a => n5151, b => n2652, outb => n2700);
   U3823 : xor2 port map( a => n5152, b => n2655, outb => n364);
   U3824 : xor2 port map( a => n5153, b => n2661, outb => n2706);
   U3825 : xor2 port map( a => n5154, b => n2663, outb => n2709);
   U3826 : xor2 port map( a => n5155, b => n2666, outb => n2712);
   U3827 : xor2 port map( a => n5156, b => n2669, outb => n2715);
   U3828 : xor2 port map( a => n5157, b => n2673, outb => n2721);
   U3829 : xor2 port map( a => n5158, b => n2675, outb => n2724);
   U3830 : xor2 port map( a => n5159, b => n2678, outb => n2727);
   U3831 : xor2 port map( a => n5160, b => n2681, outb => n2730);
   U3832 : xor2 port map( a => n5161, b => n2684, outb => n2733);
   U3833 : xor2 port map( a => n5162, b => n2687, outb => n2736);
   U3834 : xor2 port map( a => n5163, b => n2690, outb => n2739);
   U3835 : xor2 port map( a => n5164, b => n2693, outb => n2741);
   U3836 : xor2 port map( a => n5165, b => n2696, outb => n368);
   U3837 : xor2 port map( a => n5166, b => n2702, outb => n2747);
   U3838 : xor2 port map( a => n5167, b => n2704, outb => n2750);
   U3839 : xor2 port map( a => n5168, b => n2707, outb => n2753);
   U3840 : xor2 port map( a => n5169, b => n2710, outb => n2756);
   U3841 : xor2 port map( a => n5170, b => n2713, outb => n2759);
   U3842 : xor2 port map( a => n5171, b => n2717, outb => n2765);
   U3843 : xor2 port map( a => n5172, b => n2719, outb => n2768);
   U3844 : xor2 port map( a => n5173, b => n2722, outb => n2771);
   U3845 : xor2 port map( a => n5174, b => n2725, outb => n2774);
   U3846 : xor2 port map( a => n5175, b => n2728, outb => n2777);
   U3847 : xor2 port map( a => n5176, b => n2731, outb => n2780);
   U3848 : xor2 port map( a => n5177, b => n2734, outb => n2782);
   U3849 : xor2 port map( a => n5178, b => n2737, outb => n372);
   U3850 : xor2 port map( a => n5179, b => n2743, outb => n2788);
   U3851 : xor2 port map( a => n5180, b => n2745, outb => n2791);
   U3852 : xor2 port map( a => n5181, b => n2748, outb => n2794);
   U3853 : xor2 port map( a => n5182, b => n2751, outb => n2797);
   U3854 : xor2 port map( a => n5183, b => n2754, outb => n2800);
   U3855 : xor2 port map( a => n5184, b => n2757, outb => n2803);
   U3856 : xor2 port map( a => n5185, b => n2761, outb => n2809);
   U3857 : xor2 port map( a => n5186, b => n2763, outb => n2812);
   U3858 : xor2 port map( a => n5187, b => n2766, outb => n2815);
   U3859 : xor2 port map( a => n5188, b => n2769, outb => n2818);
   U3860 : xor2 port map( a => n5189, b => n2772, outb => n2821);
   U3861 : xor2 port map( a => n5190, b => n2775, outb => n2824);
   U3862 : xor2 port map( a => n5191, b => n2778, outb => n377);
   U3863 : xor2 port map( a => n5192, b => n2784, outb => n4158);
   U3864 : xor2 port map( a => n5193, b => n2786, outb => n4162);
   U3865 : xor2 port map( a => n5194, b => n2789, outb => n4166);
   U3866 : xor2 port map( a => n5195, b => n2792, outb => n4170);
   U3867 : xor2 port map( a => n5196, b => n2795, outb => n4174);
   U3868 : xor2 port map( a => n5197, b => n2798, outb => n4178);
   U3869 : inv port map( inb => n2822, outb => n5090);
   U3870 : xor2 port map( a => n5198, b => n2801, outb => n379);
   U3871 : xor2 port map( a => n5199, b => n2822, outb => n383);
   U3872 : xor2 port map( a => n3894, b => mult_125_G3_ab_2_14_port, outb => 
                           n2539);
   U3873 : xor2 port map( a => n3895, b => n3896, outb => n5108);
   U3874 : xor2 port map( a => n3897, b => n3898, outb => n5109);
   U3875 : xor2 port map( a => n3899, b => n3900, outb => n5110);
   U3876 : xor2 port map( a => n3901, b => n3902, outb => n5111);
   U3877 : xor2 port map( a => n3903, b => n3904, outb => n5112);
   U3878 : xor2 port map( a => mult_125_G3_ab_13_15_port, b => 
                           mult_125_G3_ab_14_14_port, outb => n5113);
   U3879 : xor2 port map( a => n3905, b => n837, outb => n2542);
   U3880 : xor2 port map( a => mult_125_G3_ab_3_13_port, b => n841, outb => 
                           n5114);
   U3881 : xor2 port map( a => mult_125_G3_ab_4_13_port, b => n843, outb => 
                           n2544);
   U3882 : xor2 port map( a => mult_125_G3_ab_5_13_port, b => n845, outb => 
                           n2547);
   U3883 : xor2 port map( a => mult_125_G3_ab_6_13_port, b => n847, outb => 
                           n2550);
   U3884 : xor2 port map( a => n3912, b => n3910, outb => n2553);
   U3885 : xor2 port map( a => mult_125_G3_ab_8_13_port, b => n851, outb => 
                           n2556);
   U3886 : xor2 port map( a => n3915, b => n3913, outb => n2559);
   U3887 : xor2 port map( a => mult_125_G3_ab_10_13_port, b => n855, outb => 
                           n2562);
   U3888 : xor2 port map( a => n3918, b => n3916, outb => n2565);
   U3889 : xor2 port map( a => mult_125_G3_ab_12_13_port, b => n859, outb => 
                           n2568);
   U3890 : xor2 port map( a => n3921, b => n3919, outb => n2571);
   U3891 : xor2 port map( a => mult_125_G3_ab_14_13_port, b => n863, outb => 
                           n2574);
   U3892 : xor2 port map( a => mult_125_G3_ab_15_13_port, b => n3922, outb => 
                           n2576);
   U3893 : xor2 port map( a => n868, b => mult_125_G3_ab_2_12_port, outb => 
                           n2580);
   U3894 : xor2 port map( a => n3926, b => n3924, outb => n5115);
   U3895 : xor2 port map( a => mult_125_G3_ab_4_12_port, b => n872, outb => 
                           n2582);
   U3896 : xor2 port map( a => mult_125_G3_ab_5_12_port, b => n3927, outb => 
                           n5116);
   U3897 : xor2 port map( a => n3931, b => n3929, outb => n5117);
   U3898 : xor2 port map( a => mult_125_G3_ab_7_12_port, b => n878, outb => 
                           n5118);
   U3899 : xor2 port map( a => n3934, b => n3932, outb => n5119);
   U3900 : xor2 port map( a => mult_125_G3_ab_9_12_port, b => n882, outb => 
                           n5120);
   U3901 : xor2 port map( a => n3937, b => n3935, outb => n5121);
   U3902 : xor2 port map( a => mult_125_G3_ab_11_12_port, b => n886, outb => 
                           n5122);
   U3903 : xor2 port map( a => n3940, b => n3938, outb => n5123);
   U3904 : xor2 port map( a => mult_125_G3_ab_13_12_port, b => n890, outb => 
                           n5124);
   U3905 : xor2 port map( a => n3943, b => n3941, outb => n5125);
   U3906 : xor2 port map( a => n5200, b => n894, outb => n5126);
   U3907 : xor2 port map( a => n897, b => mult_125_G3_ab_2_11_port, outb => 
                           n2586);
   U3908 : xor2 port map( a => mult_125_G3_ab_3_11_port, b => n900, outb => 
                           n5127);
   U3909 : xor2 port map( a => n3947, b => n3946, outb => n2588);
   U3910 : xor2 port map( a => mult_125_G3_ab_5_11_port, b => n904, outb => 
                           n5128);
   U3911 : xor2 port map( a => mult_125_G3_ab_6_11_port, b => n906, outb => 
                           n2591);
   U3912 : xor2 port map( a => n3952, b => n3951, outb => n2594);
   U3913 : xor2 port map( a => mult_125_G3_ab_8_11_port, b => n910, outb => 
                           n2597);
   U3914 : xor2 port map( a => n3955, b => n3953, outb => n2600);
   U3915 : xor2 port map( a => mult_125_G3_ab_10_11_port, b => n914, outb => 
                           n2603);
   U3916 : xor2 port map( a => n3958, b => n3956, outb => n2606);
   U3917 : xor2 port map( a => mult_125_G3_ab_12_11_port, b => n918, outb => 
                           n2609);
   U3918 : xor2 port map( a => n3961, b => n3959, outb => n2612);
   U3919 : xor2 port map( a => mult_125_G3_ab_14_11_port, b => n922, outb => 
                           n2615);
   U3920 : xor2 port map( a => n924, b => n925, outb => n2617);
   U3921 : xor2 port map( a => n928, b => mult_125_G3_ab_2_10_port, outb => 
                           n2621);
   U3922 : xor2 port map( a => n3965, b => n3963, outb => n5129);
   U3923 : xor2 port map( a => mult_125_G3_ab_4_10_port, b => n932, outb => 
                           n2623);
   U3924 : xor2 port map( a => n934, b => n935, outb => n5130);
   U3925 : xor2 port map( a => mult_125_G3_ab_6_10_port, b => n937, outb => 
                           n2626);
   U3926 : xor2 port map( a => mult_125_G3_ab_7_10_port, b => n939, outb => 
                           n5131);
   U3927 : xor2 port map( a => n3971, b => n3972, outb => n5132);
   U3928 : xor2 port map( a => mult_125_G3_ab_9_10_port, b => n943, outb => 
                           n5133);
   U3929 : xor2 port map( a => n3975, b => n3973, outb => n5134);
   U3930 : xor2 port map( a => mult_125_G3_ab_11_10_port, b => n947, outb => 
                           n5135);
   U3931 : xor2 port map( a => n3978, b => n3976, outb => n5136);
   U3932 : xor2 port map( a => mult_125_G3_ab_13_10_port, b => n951, outb => 
                           n5137);
   U3933 : xor2 port map( a => n3981, b => n3979, outb => n5138);
   U3934 : xor2 port map( a => n5201, b => n955, outb => n5139);
   U3935 : xor2 port map( a => n958, b => mult_125_G3_ab_2_9_port, outb => 
                           n2630);
   U3936 : xor2 port map( a => n3984, b => n3982, outb => n5140);
   U3937 : xor2 port map( a => mult_125_G3_ab_4_9_port, b => n962, outb => 
                           n2632);
   U3938 : xor2 port map( a => mult_125_G3_ab_5_9_port, b => n964, outb => 
                           n5141);
   U3939 : xor2 port map( a => mult_125_G3_ab_6_9_port, b => n966, outb => 
                           n2635);
   U3940 : xor2 port map( a => mult_125_G3_ab_7_9_port, b => n968, outb => 
                           n5142);
   U3941 : xor2 port map( a => n3992, b => n3990, outb => n2638);
   U3942 : xor2 port map( a => n3994, b => n3993, outb => n2641);
   U3943 : xor2 port map( a => mult_125_G3_ab_10_9_port, b => n974, outb => 
                           n2644);
   U3944 : xor2 port map( a => n3997, b => n3995, outb => n2647);
   U3945 : xor2 port map( a => mult_125_G3_ab_12_9_port, b => n978, outb => 
                           n2650);
   U3946 : xor2 port map( a => n4000, b => n3998, outb => n2653);
   U3947 : xor2 port map( a => mult_125_G3_ab_14_9_port, b => n982, outb => 
                           n2656);
   U3948 : xor2 port map( a => n984, b => n985, outb => n2658);
   U3949 : xor2 port map( a => n988, b => mult_125_G3_ab_2_8_port, outb => 
                           n2662);
   U3950 : xor2 port map( a => n4004, b => n4002, outb => n5143);
   U3951 : xor2 port map( a => n4006, b => n992, outb => n2664);
   U3952 : xor2 port map( a => n4008, b => n4007, outb => n5144);
   U3953 : xor2 port map( a => mult_125_G3_ab_6_8_port, b => n996, outb => 
                           n2667);
   U3954 : xor2 port map( a => n4011, b => n4009, outb => n5145);
   U3955 : xor2 port map( a => mult_125_G3_ab_8_8_port, b => n1000, outb => 
                           n2670);
   U3956 : xor2 port map( a => mult_125_G3_ab_9_8_port, b => n1002, outb => 
                           n5146);
   U3957 : xor2 port map( a => n4015, b => n4016, outb => n5147);
   U3958 : xor2 port map( a => mult_125_G3_ab_11_8_port, b => n1006, outb => 
                           n5148);
   U3959 : xor2 port map( a => n4019, b => n4017, outb => n5149);
   U3960 : xor2 port map( a => mult_125_G3_ab_13_8_port, b => n1010, outb => 
                           n5150);
   U3961 : xor2 port map( a => n4022, b => n4020, outb => n5151);
   U3962 : xor2 port map( a => n5202, b => n1014, outb => n5152);
   U3963 : xor2 port map( a => n1017, b => mult_125_G3_ab_2_7_port, outb => 
                           n2674);
   U3964 : xor2 port map( a => mult_125_G3_ab_3_7_port, b => n1020, outb => 
                           n5153);
   U3965 : xor2 port map( a => n4026, b => n4025, outb => n2676);
   U3966 : xor2 port map( a => mult_125_G3_ab_5_7_port, b => n1024, outb => 
                           n5154);
   U3967 : xor2 port map( a => n4029, b => n4027, outb => n2679);
   U3968 : xor2 port map( a => mult_125_G3_ab_7_7_port, b => n1028, outb => 
                           n5155);
   U3969 : xor2 port map( a => n4032, b => n4030, outb => n2682);
   U3970 : xor2 port map( a => mult_125_G3_ab_9_7_port, b => n1032, outb => 
                           n5156);
   U3971 : xor2 port map( a => n4035, b => n4033, outb => n2685);
   U3972 : xor2 port map( a => n4037, b => n4036, outb => n2688);
   U3973 : xor2 port map( a => mult_125_G3_ab_12_7_port, b => n1038, outb => 
                           n2691);
   U3974 : xor2 port map( a => n4040, b => n4038, outb => n2694);
   U3975 : xor2 port map( a => mult_125_G3_ab_14_7_port, b => n1042, outb => 
                           n2697);
   U3976 : xor2 port map( a => n1044, b => n1045, outb => n2699);
   U3977 : xor2 port map( a => n1048, b => mult_125_G3_ab_2_6_port, outb => 
                           n2703);
   U3978 : xor2 port map( a => n4044, b => n4042, outb => n5157);
   U3979 : xor2 port map( a => mult_125_G3_ab_4_6_port, b => n1052, outb => 
                           n2705);
   U3980 : xor2 port map( a => n1054, b => n1055, outb => n5158);
   U3981 : xor2 port map( a => mult_125_G3_ab_6_6_port, b => n1057, outb => 
                           n2708);
   U3982 : xor2 port map( a => n4049, b => n4047, outb => n5159);
   U3983 : xor2 port map( a => mult_125_G3_ab_8_6_port, b => n1061, outb => 
                           n2711);
   U3984 : xor2 port map( a => n1063, b => n1064, outb => n5160);
   U3985 : xor2 port map( a => mult_125_G3_ab_10_6_port, b => n1066, outb => 
                           n2714);
   U3986 : xor2 port map( a => mult_125_G3_ab_11_6_port, b => n1068, outb => 
                           n5161);
   U3987 : xor2 port map( a => n4055, b => n4056, outb => n5162);
   U3988 : xor2 port map( a => mult_125_G3_ab_13_6_port, b => n1072, outb => 
                           n5163);
   U3989 : xor2 port map( a => n4059, b => n4057, outb => n5164);
   U3990 : xor2 port map( a => n5203, b => n1076, outb => n5165);
   U3991 : xor2 port map( a => n1079, b => mult_125_G3_ab_2_5_port, outb => 
                           n2718);
   U3992 : xor2 port map( a => mult_125_G3_ab_3_5_port, b => n1082, outb => 
                           n5166);
   U3993 : xor2 port map( a => mult_125_G3_ab_4_5_port, b => n1084, outb => 
                           n2720);
   U3994 : xor2 port map( a => mult_125_G3_ab_5_5_port, b => n1086, outb => 
                           n5167);
   U3995 : xor2 port map( a => n1088, b => n1089, outb => n2723);
   U3996 : xor2 port map( a => mult_125_G3_ab_7_5_port, b => n1091, outb => 
                           n5168);
   U3997 : xor2 port map( a => mult_125_G3_ab_8_5_port, b => n1093, outb => 
                           n2726);
   U3998 : xor2 port map( a => mult_125_G3_ab_9_5_port, b => n1095, outb => 
                           n5169);
   U3999 : xor2 port map( a => n4071, b => n4069, outb => n2729);
   U4000 : xor2 port map( a => mult_125_G3_ab_11_5_port, b => n1099, outb => 
                           n5170);
   U4001 : xor2 port map( a => n4074, b => n4072, outb => n2732);
   U4002 : xor2 port map( a => n4076, b => n1103, outb => n2735);
   U4003 : xor2 port map( a => mult_125_G3_ab_14_5_port, b => n1105, outb => 
                           n2738);
   U4004 : xor2 port map( a => n1107, b => n1108, outb => n2740);
   U4005 : xor2 port map( a => n1111, b => mult_125_G3_ab_2_4_port, outb => 
                           n2744);
   U4006 : xor2 port map( a => n4080, b => n4078, outb => n5171);
   U4007 : xor2 port map( a => mult_125_G3_ab_4_4_port, b => n1115, outb => 
                           n2746);
   U4008 : xor2 port map( a => n1117, b => n1118, outb => n5172);
   U4009 : xor2 port map( a => mult_125_G3_ab_6_4_port, b => n1120, outb => 
                           n2749);
   U4010 : xor2 port map( a => n1122, b => n1123, outb => n5173);
   U4011 : xor2 port map( a => mult_125_G3_ab_8_4_port, b => n1125, outb => 
                           n2752);
   U4012 : xor2 port map( a => mult_125_G3_ab_9_4_port, b => n1127, outb => 
                           n5174);
   U4013 : xor2 port map( a => mult_125_G3_ab_10_4_port, b => n1129, outb => 
                           n2755);
   U4014 : xor2 port map( a => n1131, b => n1132, outb => n5175);
   U4015 : xor2 port map( a => mult_125_G3_ab_12_4_port, b => n1134, outb => 
                           n2758);
   U4016 : xor2 port map( a => mult_125_G3_ab_13_4_port, b => n1136, outb => 
                           n5176);
   U4017 : xor2 port map( a => mult_125_G3_ab_14_4_port, b => n1138, outb => 
                           n5177);
   U4018 : xor2 port map( a => mult_125_G3_ab_15_4_port, b => n1141, outb => 
                           n5178);
   U4019 : xor2 port map( a => n1144, b => mult_125_G3_ab_2_3_port, outb => 
                           n2762);
   U4020 : xor2 port map( a => mult_125_G3_ab_3_3_port, b => n1147, outb => 
                           n5179);
   U4021 : xor2 port map( a => mult_125_G3_ab_4_3_port, b => n1149, outb => 
                           n2764);
   U4022 : xor2 port map( a => mult_125_G3_ab_5_3_port, b => n1151, outb => 
                           n5180);
   U4023 : xor2 port map( a => mult_125_G3_ab_6_3_port, b => n1153, outb => 
                           n2767);
   U4024 : xor2 port map( a => mult_125_G3_ab_7_3_port, b => n1155, outb => 
                           n5181);
   U4025 : xor2 port map( a => mult_125_G3_ab_8_3_port, b => n1157, outb => 
                           n2770);
   U4026 : xor2 port map( a => mult_125_G3_ab_9_3_port, b => n1159, outb => 
                           n5182);
   U4027 : xor2 port map( a => mult_125_G3_ab_10_3_port, b => n1161, outb => 
                           n2773);
   U4028 : xor2 port map( a => mult_125_G3_ab_11_3_port, b => n1163, outb => 
                           n5183);
   U4029 : xor2 port map( a => n4109, b => n4107, outb => n2776);
   U4030 : xor2 port map( a => mult_125_G3_ab_13_3_port, b => n1167, outb => 
                           n5184);
   U4031 : xor2 port map( a => mult_125_G3_ab_14_3_port, b => n1169, outb => 
                           n2779);
   U4032 : xor2 port map( a => mult_125_G3_ab_15_3_port, b => n1171, outb => 
                           n2781);
   U4033 : xor2 port map( a => n1174, b => mult_125_G3_ab_2_2_port, outb => 
                           n2785);
   U4034 : xor2 port map( a => n4115, b => n4113, outb => n5185);
   U4035 : xor2 port map( a => mult_125_G3_ab_4_2_port, b => n1178, outb => 
                           n2787);
   U4036 : xor2 port map( a => mult_125_G3_ab_5_2_port, b => n1180, outb => 
                           n5186);
   U4037 : xor2 port map( a => mult_125_G3_ab_6_2_port, b => n1182, outb => 
                           n2790);
   U4038 : xor2 port map( a => n1184, b => n1185, outb => n5187);
   U4039 : xor2 port map( a => mult_125_G3_ab_8_2_port, b => n1187, outb => 
                           n2793);
   U4040 : xor2 port map( a => mult_125_G3_ab_9_2_port, b => n1189, outb => 
                           n5188);
   U4041 : xor2 port map( a => mult_125_G3_ab_10_2_port, b => n1191, outb => 
                           n2796);
   U4042 : xor2 port map( a => mult_125_G3_ab_11_2_port, b => n1193, outb => 
                           n5189);
   U4043 : xor2 port map( a => mult_125_G3_ab_12_2_port, b => n1195, outb => 
                           n2799);
   U4044 : xor2 port map( a => mult_125_G3_ab_13_2_port, b => n1197, outb => 
                           n5190);
   U4045 : xor2 port map( a => mult_125_G3_ab_14_2_port, b => n1199, outb => 
                           n2802);
   U4046 : xor2 port map( a => n5087, b => n4130, outb => n5191);
   U4047 : xor2 port map( a => n4133, b => mult_125_G3_ab_2_1_port, outb => 
                           n2806);
   U4048 : xor2 port map( a => n4134, b => n4132, outb => n5192);
   U4049 : xor2 port map( a => mult_125_G3_ab_4_1_port, b => n4136, outb => 
                           n2808);
   U4050 : xor2 port map( a => mult_125_G3_ab_5_1_port, b => n1210, outb => 
                           n5204);
   U4051 : xor2 port map( a => n4139, b => n1212, outb => n2811);
   U4052 : xor2 port map( a => n5205, b => n1214, outb => n5194);
   U4053 : xor2 port map( a => mult_125_G3_ab_8_1_port, b => n4140, outb => 
                           n2814);
   U4054 : xor2 port map( a => n5206, b => n1218, outb => n5195);
   U4055 : xor2 port map( a => n4145, b => n1220, outb => n2817);
   U4056 : xor2 port map( a => n5207, b => n1222, outb => n5196);
   U4057 : xor2 port map( a => n4148, b => n1224, outb => n2820);
   U4058 : xor2 port map( a => n5208, b => n1226, outb => n5197);
   U4059 : xor2 port map( a => n4151, b => n4149, outb => n2823);
   U4060 : xor2 port map( a => n5209, b => n1230, outb => n5198);
   U4061 : xor2 port map( a => mult_125_G3_ab_15_0_port, b => n1258, outb => 
                           n5199);
   U4062 : xor2 port map( a => mult_125_G3_ab_11_0_port, b => n1250, outb => 
                           n2825);
   U4063 : xor2 port map( a => mult_125_G3_ab_9_0_port, b => n1246, outb => 
                           n2826);
   U4064 : xor2 port map( a => mult_125_G3_ab_7_0_port, b => n1242, outb => 
                           n2827);
   U4065 : xor2 port map( a => mult_125_G3_ab_5_0_port, b => n1238, outb => 
                           n2828);
   U4066 : xor2 port map( a => mult_125_G3_ab_3_0_port, b => n1234, outb => 
                           n2829);
   U4067 : xor2 port map( a => n380, b => mult_125_G3_ZA, outb => n2830);
   U4068 : xor2 port map( a => mult_125_G3_ab_13_0_port, b => n1254, outb => 
                           n2831);
   U4069 : xor2 port map( a => n4774, b => adder_mem_array_3_26_port, outb => 
                           n3429);
   U4070 : xor2 port map( a => n4772, b => adder_mem_array_3_24_port, outb => 
                           n3433);
   U4071 : xor2 port map( a => n4770, b => adder_mem_array_3_22_port, outb => 
                           n3437);
   U4072 : xor2 port map( a => n4768, b => adder_mem_array_3_20_port, outb => 
                           n3441);
   U4073 : xor2 port map( a => n4766, b => adder_mem_array_3_18_port, outb => 
                           n3445);
   U4074 : xor2 port map( a => n4764, b => adder_mem_array_3_16_port, outb => 
                           n3452);
   U4075 : xor2 port map( a => n4762, b => adder_mem_array_3_14_port, outb => 
                           n3456);
   U4076 : xor2 port map( a => n4760, b => adder_mem_array_3_12_port, outb => 
                           n3460);
   U4077 : xor2 port map( a => n4758, b => adder_mem_array_3_10_port, outb => 
                           n3464);
   U4078 : xor2 port map( a => n4756, b => adder_mem_array_3_8_port, outb => 
                           n3468);
   U4079 : xor2 port map( a => n4754, b => adder_mem_array_3_6_port, outb => 
                           n3474);
   U4080 : xor2 port map( a => n4752, b => adder_mem_array_3_4_port, outb => 
                           n3478);
   U4081 : xor2 port map( a => n4750, b => adder_mem_array_3_2_port, outb => 
                           n3482);
   U4082 : xor2 port map( a => n5107, b => adder_mem_array_3_32_port, outb => 
                           n3599);
   U4083 : xor2 port map( a => n4840, b => adder_mem_array_3_30_port, outb => 
                           n3601);
   U4084 : xor2 port map( a => n4838, b => adder_mem_array_3_28_port, outb => 
                           n3605);
   U4085 : oai22 port map( a => n5211, b => n5212, c => n1260, d => n4179, outb
                           => n5210);
   U4086 : aoi22 port map( a => mult_125_G2_ab_2_15_port, b => 
                           mult_125_G2_ab_3_14_port, c => n5210, d => n5214, 
                           outb => n5213);
   U4087 : oai22 port map( a => n4180, b => n4181, c => n5213, d => n1262, outb
                           => n5215);
   U4088 : aoi22 port map( a => mult_125_G2_ab_4_15_port, b => 
                           mult_125_G2_ab_5_14_port, c => n5215, d => n5217, 
                           outb => n5216);
   U4089 : oai22 port map( a => n4182, b => n4183, c => n5216, d => n1264, outb
                           => n5218);
   U4090 : aoi22 port map( a => mult_125_G2_ab_6_15_port, b => 
                           mult_125_G2_ab_7_14_port, c => n5218, d => n5220, 
                           outb => n5219);
   U4091 : oai22 port map( a => n4184, b => n4185, c => n5219, d => n1266, outb
                           => n5221);
   U4092 : aoi22 port map( a => mult_125_G2_ab_8_15_port, b => 
                           mult_125_G2_ab_9_14_port, c => n5221, d => n5223, 
                           outb => n5222);
   U4093 : oai22 port map( a => n4186, b => n4187, c => n5222, d => n1268, outb
                           => n5224);
   U4094 : aoi22 port map( a => mult_125_G2_ab_10_15_port, b => 
                           mult_125_G2_ab_11_14_port, c => n5224, d => n5226, 
                           outb => n5225);
   U4095 : oai22 port map( a => n4188, b => n4189, c => n5225, d => n1270, outb
                           => n5227);
   U4096 : aoi22 port map( a => mult_125_G2_ab_12_15_port, b => 
                           mult_125_G2_ab_13_14_port, c => n5227, d => n5229, 
                           outb => n5228);
   U4097 : aoi22 port map( a => mult_125_G2_ab_13_15_port, b => 
                           mult_125_G2_ab_14_14_port, c => n5231, d => n5232, 
                           outb => n5230);
   U4098 : aoi22 port map( a => mult_125_G2_ab_14_15_port, b => 
                           mult_125_G2_ab_15_14_port, c => n5233, d => n5234, 
                           outb => n313);
   U4099 : inv port map( inb => n4207, outb => n1303);
   U4100 : aoi22 port map( a => n1303, b => mult_125_G2_ab_15_13_port, c => 
                           n5235, d => n2874, outb => n315);
   U4101 : aoi22 port map( a => n1332, b => mult_125_G2_ab_15_12_port, c => 
                           n5236, d => n2870, outb => n317);
   U4102 : oai22 port map( a => n1363, b => n1362, c => n5238, d => n2915, outb
                           => n5237);
   U4103 : inv port map( inb => n1379, outb => n4257);
   U4104 : aoi22 port map( a => n1393, b => mult_125_G2_ab_15_10_port, c => 
                           n5239, d => n2911, outb => n321);
   U4105 : oai22 port map( a => n1423, b => n1422, c => n5241, d => n2956, outb
                           => n5240);
   U4106 : inv port map( inb => n1442, outb => n4301);
   U4107 : aoi22 port map( a => n1452, b => mult_125_G2_ab_15_8_port, c => 
                           n5242, d => n2952, outb => n325);
   U4108 : oai22 port map( a => n1483, b => n1482, c => n5244, d => n2997, outb
                           => n5243);
   U4109 : inv port map( inb => n1508, outb => n4341);
   U4110 : aoi22 port map( a => n1514, b => mult_125_G2_ab_15_6_port, c => 
                           n5245, d => n2993, outb => n329);
   U4111 : oai22 port map( a => n1546, b => n1545, c => n5247, d => n3038, outb
                           => n5246);
   U4112 : aoi22 port map( a => n5248, b => mult_125_G2_ab_15_4_port, c => 
                           n1577, d => n3034, outb => n333);
   U4113 : aoi22 port map( a => n1609, b => mult_125_G2_ab_15_3_port, c => 
                           n5249, d => n3079, outb => n335);
   U4114 : oai22 port map( a => n4415, b => n5250, c => n1638, d => n3075, outb
                           => n338);
   U4115 : aoi22 port map( a => n1668, b => mult_125_G2_ab_15_1_port, c => 
                           n5251, d => n3098, outb => n340);
   U4116 : aoi22 port map( a => n1696, b => mult_125_G2_ab_15_0_port, c => 
                           n5252, d => n5253, outb => n342);
   U4117 : aoi22 port map( a => adder_mem_array_2_1_port, b => n2167, c => 
                           n5254, d => n3484, outb => n3544);
   U4118 : oai22 port map( a => n4780, b => n4781, c => n3544, d => n2168, outb
                           => n3541);
   U4119 : aoi22 port map( a => multiplier_sigs_1_3_port, b => 
                           adder_mem_array_2_3_port, c => n3541, d => n5255, 
                           outb => n3540);
   U4120 : oai22 port map( a => n4782, b => n4783, c => n3540, d => n2170, outb
                           => n3537);
   U4121 : aoi22 port map( a => multiplier_sigs_1_5_port, b => 
                           adder_mem_array_2_5_port, c => n3537, d => n5256, 
                           outb => n3536);
   U4122 : oai22 port map( a => n4784, b => n4785, c => n3536, d => n2172, outb
                           => n3533);
   U4123 : aoi22 port map( a => multiplier_sigs_1_7_port, b => 
                           adder_mem_array_2_7_port, c => n3533, d => n5257, 
                           outb => n3532);
   U4124 : oai22 port map( a => n4786, b => n4787, c => n3532, d => n2174, outb
                           => n3529);
   U4125 : aoi22 port map( a => multiplier_sigs_1_9_port, b => 
                           adder_mem_array_2_9_port, c => n3529, d => n5258, 
                           outb => n3528);
   U4126 : oai22 port map( a => n4788, b => n4789, c => n3528, d => n2176, outb
                           => n3525);
   U4127 : aoi22 port map( a => multiplier_sigs_1_11_port, b => 
                           adder_mem_array_2_11_port, c => n3525, d => n5259, 
                           outb => n3524);
   U4128 : oai22 port map( a => n4790, b => n4791, c => n3524, d => n2178, outb
                           => n3521);
   U4129 : aoi22 port map( a => multiplier_sigs_1_13_port, b => 
                           adder_mem_array_2_13_port, c => n3521, d => n5260, 
                           outb => n3520);
   U4130 : oai22 port map( a => n4792, b => n4793, c => n3520, d => n2180, outb
                           => n3517);
   U4131 : aoi22 port map( a => multiplier_sigs_1_15_port, b => 
                           adder_mem_array_2_15_port, c => n3517, d => n5261, 
                           outb => n3516);
   U4132 : oai22 port map( a => n4794, b => n4795, c => n3516, d => n2182, outb
                           => n3513);
   U4133 : aoi22 port map( a => multiplier_sigs_1_17_port, b => 
                           adder_mem_array_2_17_port, c => n3513, d => n5262, 
                           outb => n3512);
   U4134 : oai22 port map( a => n4796, b => n4797, c => n3512, d => n2184, outb
                           => n3509);
   U4135 : aoi22 port map( a => multiplier_sigs_1_19_port, b => 
                           adder_mem_array_2_19_port, c => n3509, d => n5263, 
                           outb => n3508);
   U4136 : oai22 port map( a => n4798, b => n4799, c => n3508, d => n2186, outb
                           => n3505);
   U4137 : aoi22 port map( a => multiplier_sigs_1_21_port, b => 
                           adder_mem_array_2_21_port, c => n3505, d => n5264, 
                           outb => n3504);
   U4138 : oai22 port map( a => n4800, b => n4801, c => n3504, d => n2188, outb
                           => n3501);
   U4139 : aoi22 port map( a => multiplier_sigs_1_23_port, b => 
                           adder_mem_array_2_23_port, c => n3501, d => n5265, 
                           outb => n3500);
   U4140 : oai22 port map( a => n4802, b => n4803, c => n3500, d => n2190, outb
                           => n3497);
   U4141 : aoi22 port map( a => multiplier_sigs_1_25_port, b => 
                           adder_mem_array_2_25_port, c => n3497, d => n5266, 
                           outb => n3496);
   U4142 : oai22 port map( a => n4804, b => n4805, c => n3496, d => n2192, outb
                           => n3493);
   U4143 : aoi22 port map( a => multiplier_sigs_1_27_port, b => 
                           adder_mem_array_2_27_port, c => n3493, d => n5267, 
                           outb => n3492);
   U4144 : oai22 port map( a => n4806, b => n4807, c => n3492, d => n2194, outb
                           => n3489);
   U4145 : aoi22 port map( a => multiplier_sigs_1_29_port, b => 
                           adder_mem_array_2_29_port, c => n3489, d => n5268, 
                           outb => n3488);
   U4146 : oai22 port map( a => n4808, b => n4809, c => n3488, d => n2196, outb
                           => n2199);
   U4147 : nand2 port map( a => n5269, b => n5270, outb => n2198);
   U4148 : xor2 port map( a => n5210, b => n4887, outb => n2842);
   U4149 : xor2 port map( a => n5271, b => n5213, outb => n2845);
   U4150 : xor2 port map( a => n5215, b => n4888, outb => n2848);
   U4151 : xor2 port map( a => n5272, b => n5216, outb => n2851);
   U4152 : xor2 port map( a => n5218, b => n4889, outb => n2854);
   U4153 : xor2 port map( a => n5273, b => n5219, outb => n2857);
   U4154 : xor2 port map( a => n5221, b => n4890, outb => n2860);
   U4155 : xor2 port map( a => n5274, b => n5222, outb => n2863);
   U4156 : xor2 port map( a => n5224, b => n4891, outb => n2866);
   U4157 : xor2 port map( a => n5275, b => n5225, outb => n2869);
   U4158 : xor2 port map( a => n5227, b => n4892, outb => n2872);
   U4159 : xor2 port map( a => n5276, b => n5231, outb => n2874);
   U4160 : xor2 port map( a => n5230, b => n4893, outb => n316);
   U4161 : xor2 port map( a => n5277, b => n2835, outb => n2880);
   U4162 : xor2 port map( a => n5278, b => n2838, outb => n2886);
   U4163 : xor2 port map( a => n5279, b => n2840, outb => n2889);
   U4164 : xor2 port map( a => n5280, b => n2843, outb => n2892);
   U4165 : xor2 port map( a => n5281, b => n2846, outb => n2895);
   U4166 : xor2 port map( a => n5282, b => n2849, outb => n2898);
   U4167 : xor2 port map( a => n5283, b => n2852, outb => n2901);
   U4168 : xor2 port map( a => n5284, b => n2855, outb => n2904);
   U4169 : xor2 port map( a => n5285, b => n2858, outb => n2907);
   U4170 : xor2 port map( a => n5286, b => n2861, outb => n2910);
   U4171 : xor2 port map( a => n5287, b => n2864, outb => n2913);
   U4172 : xor2 port map( a => n5288, b => n2867, outb => n2915);
   U4173 : xor2 port map( a => n5289, b => n2870, outb => n320);
   U4174 : xor2 port map( a => n5290, b => n2876, outb => n2921);
   U4175 : xor2 port map( a => n5291, b => n2878, outb => n2924);
   U4176 : xor2 port map( a => n5292, b => n2882, outb => n2930);
   U4177 : xor2 port map( a => n5293, b => n2884, outb => n2933);
   U4178 : xor2 port map( a => n5294, b => n2887, outb => n2936);
   U4179 : xor2 port map( a => n5295, b => n2890, outb => n2939);
   U4180 : xor2 port map( a => n5296, b => n2893, outb => n2942);
   U4181 : xor2 port map( a => n5297, b => n2896, outb => n2945);
   U4182 : xor2 port map( a => n5298, b => n2899, outb => n2948);
   U4183 : xor2 port map( a => n5299, b => n2902, outb => n2951);
   U4184 : xor2 port map( a => n5300, b => n2905, outb => n2954);
   U4185 : xor2 port map( a => n5301, b => n2908, outb => n2956);
   U4186 : xor2 port map( a => n5302, b => n2911, outb => n324);
   U4187 : xor2 port map( a => n5303, b => n2917, outb => n2962);
   U4188 : xor2 port map( a => n5304, b => n2919, outb => n2965);
   U4189 : xor2 port map( a => n5305, b => n2922, outb => n2968);
   U4190 : xor2 port map( a => n5306, b => n2926, outb => n2974);
   U4191 : xor2 port map( a => n5307, b => n2928, outb => n2977);
   U4192 : xor2 port map( a => n5308, b => n2931, outb => n2980);
   U4193 : xor2 port map( a => n5309, b => n2934, outb => n2983);
   U4194 : xor2 port map( a => n5310, b => n2937, outb => n2986);
   U4195 : xor2 port map( a => n5311, b => n2940, outb => n2989);
   U4196 : xor2 port map( a => n5312, b => n2943, outb => n2992);
   U4197 : xor2 port map( a => n5313, b => n2946, outb => n2995);
   U4198 : xor2 port map( a => n5314, b => n2949, outb => n2997);
   U4199 : xor2 port map( a => n5315, b => n2952, outb => n328);
   U4200 : xor2 port map( a => n5316, b => n2958, outb => n3003);
   U4201 : xor2 port map( a => n5317, b => n2960, outb => n3006);
   U4202 : xor2 port map( a => n5318, b => n2963, outb => n3009);
   U4203 : xor2 port map( a => n5319, b => n2966, outb => n3012);
   U4204 : xor2 port map( a => n5320, b => n2970, outb => n3018);
   U4205 : xor2 port map( a => n5321, b => n2972, outb => n3021);
   U4206 : xor2 port map( a => n5322, b => n2975, outb => n3024);
   U4207 : xor2 port map( a => n5323, b => n2978, outb => n3027);
   U4208 : xor2 port map( a => n5324, b => n2981, outb => n3030);
   U4209 : xor2 port map( a => n5325, b => n2984, outb => n3033);
   U4210 : xor2 port map( a => n5326, b => n2987, outb => n3036);
   U4211 : xor2 port map( a => n5327, b => n2990, outb => n3038);
   U4212 : xor2 port map( a => n5328, b => n2993, outb => n332);
   U4213 : xor2 port map( a => n5329, b => n2999, outb => n3044);
   U4214 : xor2 port map( a => n5330, b => n3001, outb => n3047);
   U4215 : xor2 port map( a => n5331, b => n3004, outb => n3050);
   U4216 : xor2 port map( a => n5332, b => n3007, outb => n3053);
   U4217 : xor2 port map( a => n5333, b => n3010, outb => n3056);
   U4218 : xor2 port map( a => n5334, b => n3014, outb => n3062);
   U4219 : xor2 port map( a => n5335, b => n3016, outb => n3065);
   U4220 : xor2 port map( a => n5336, b => n3019, outb => n3068);
   U4221 : xor2 port map( a => n5337, b => n3022, outb => n3071);
   U4222 : xor2 port map( a => n5338, b => n3025, outb => n3074);
   U4223 : xor2 port map( a => n5339, b => n3028, outb => n3077);
   U4224 : xor2 port map( a => n5340, b => n3031, outb => n3079);
   U4225 : xor2 port map( a => n5341, b => n3034, outb => n336);
   U4226 : xor2 port map( a => n5342, b => n3040, outb => n3085);
   U4227 : xor2 port map( a => n5343, b => n3042, outb => n3088);
   U4228 : xor2 port map( a => n5344, b => n3045, outb => n3091);
   U4229 : xor2 port map( a => n5345, b => n3048, outb => n3094);
   U4230 : xor2 port map( a => n5346, b => n3051, outb => n3097);
   U4231 : xor2 port map( a => n5347, b => n3054, outb => n3100);
   U4232 : xor2 port map( a => n5348, b => n3058, outb => n3106);
   U4233 : xor2 port map( a => n5349, b => n3060, outb => n3109);
   U4234 : xor2 port map( a => n5350, b => n3063, outb => n3112);
   U4235 : xor2 port map( a => n5351, b => n3066, outb => n3115);
   U4236 : xor2 port map( a => n5352, b => n3069, outb => n3118);
   U4237 : xor2 port map( a => n5353, b => n3072, outb => n3121);
   U4238 : xor2 port map( a => n5354, b => n3075, outb => n341);
   U4239 : xor2 port map( a => n5355, b => n3081, outb => n4443);
   U4240 : xor2 port map( a => n5356, b => n3083, outb => n4447);
   U4241 : xor2 port map( a => n5357, b => n3086, outb => n4451);
   U4242 : xor2 port map( a => n5358, b => n3089, outb => n4455);
   U4243 : xor2 port map( a => n5359, b => n3092, outb => n4459);
   U4244 : xor2 port map( a => n5360, b => n3095, outb => n4463);
   U4245 : inv port map( inb => n3119, outb => n5253);
   U4246 : xor2 port map( a => n5361, b => n3098, outb => n343);
   U4247 : xor2 port map( a => n5362, b => n3119, outb => n347);
   U4248 : xor2 port map( a => n4179, b => mult_125_G2_ab_2_14_port, outb => 
                           n2836);
   U4249 : xor2 port map( a => n4180, b => n4181, outb => n5271);
   U4250 : xor2 port map( a => n4182, b => n4183, outb => n5272);
   U4251 : xor2 port map( a => n4184, b => n4185, outb => n5273);
   U4252 : xor2 port map( a => n4186, b => n4187, outb => n5274);
   U4253 : xor2 port map( a => n4188, b => n4189, outb => n5275);
   U4254 : xor2 port map( a => mult_125_G2_ab_13_15_port, b => 
                           mult_125_G2_ab_14_14_port, outb => n5276);
   U4255 : xor2 port map( a => n4190, b => n1275, outb => n2839);
   U4256 : xor2 port map( a => mult_125_G2_ab_3_13_port, b => n1279, outb => 
                           n5277);
   U4257 : xor2 port map( a => mult_125_G2_ab_4_13_port, b => n1281, outb => 
                           n2841);
   U4258 : xor2 port map( a => mult_125_G2_ab_5_13_port, b => n1283, outb => 
                           n2844);
   U4259 : xor2 port map( a => mult_125_G2_ab_6_13_port, b => n1285, outb => 
                           n2847);
   U4260 : xor2 port map( a => n4197, b => n4195, outb => n2850);
   U4261 : xor2 port map( a => mult_125_G2_ab_8_13_port, b => n1289, outb => 
                           n2853);
   U4262 : xor2 port map( a => n4200, b => n4198, outb => n2856);
   U4263 : xor2 port map( a => mult_125_G2_ab_10_13_port, b => n1293, outb => 
                           n2859);
   U4264 : xor2 port map( a => n4203, b => n4201, outb => n2862);
   U4265 : xor2 port map( a => mult_125_G2_ab_12_13_port, b => n1297, outb => 
                           n2865);
   U4266 : xor2 port map( a => n4206, b => n4204, outb => n2868);
   U4267 : xor2 port map( a => mult_125_G2_ab_14_13_port, b => n1301, outb => 
                           n2871);
   U4268 : xor2 port map( a => mult_125_G2_ab_15_13_port, b => n4207, outb => 
                           n2873);
   U4269 : xor2 port map( a => n1306, b => mult_125_G2_ab_2_12_port, outb => 
                           n2877);
   U4270 : xor2 port map( a => n4211, b => n4209, outb => n5278);
   U4271 : xor2 port map( a => mult_125_G2_ab_4_12_port, b => n1310, outb => 
                           n2879);
   U4272 : xor2 port map( a => mult_125_G2_ab_5_12_port, b => n4212, outb => 
                           n5279);
   U4273 : xor2 port map( a => n4216, b => n4214, outb => n5280);
   U4274 : xor2 port map( a => mult_125_G2_ab_7_12_port, b => n1316, outb => 
                           n5281);
   U4275 : xor2 port map( a => n4219, b => n4217, outb => n5282);
   U4276 : xor2 port map( a => mult_125_G2_ab_9_12_port, b => n1320, outb => 
                           n5283);
   U4277 : xor2 port map( a => n4222, b => n4220, outb => n5284);
   U4278 : xor2 port map( a => mult_125_G2_ab_11_12_port, b => n1324, outb => 
                           n5285);
   U4279 : xor2 port map( a => n4225, b => n4223, outb => n5286);
   U4280 : xor2 port map( a => mult_125_G2_ab_13_12_port, b => n1328, outb => 
                           n5287);
   U4281 : xor2 port map( a => n4228, b => n4226, outb => n5288);
   U4282 : xor2 port map( a => n5363, b => n1332, outb => n5289);
   U4283 : xor2 port map( a => n1335, b => mult_125_G2_ab_2_11_port, outb => 
                           n2883);
   U4284 : xor2 port map( a => mult_125_G2_ab_3_11_port, b => n1338, outb => 
                           n5290);
   U4285 : xor2 port map( a => n4232, b => n4231, outb => n2885);
   U4286 : xor2 port map( a => mult_125_G2_ab_5_11_port, b => n1342, outb => 
                           n5291);
   U4287 : xor2 port map( a => mult_125_G2_ab_6_11_port, b => n1344, outb => 
                           n2888);
   U4288 : xor2 port map( a => n4237, b => n4236, outb => n2891);
   U4289 : xor2 port map( a => mult_125_G2_ab_8_11_port, b => n1348, outb => 
                           n2894);
   U4290 : xor2 port map( a => n4240, b => n4238, outb => n2897);
   U4291 : xor2 port map( a => mult_125_G2_ab_10_11_port, b => n1352, outb => 
                           n2900);
   U4292 : xor2 port map( a => n4243, b => n4241, outb => n2903);
   U4293 : xor2 port map( a => mult_125_G2_ab_12_11_port, b => n1356, outb => 
                           n2906);
   U4294 : xor2 port map( a => n4246, b => n4244, outb => n2909);
   U4295 : xor2 port map( a => mult_125_G2_ab_14_11_port, b => n1360, outb => 
                           n2912);
   U4296 : xor2 port map( a => n1362, b => n1363, outb => n2914);
   U4297 : xor2 port map( a => n1366, b => mult_125_G2_ab_2_10_port, outb => 
                           n2918);
   U4298 : xor2 port map( a => n4250, b => n4248, outb => n5292);
   U4299 : xor2 port map( a => mult_125_G2_ab_4_10_port, b => n1370, outb => 
                           n2920);
   U4300 : xor2 port map( a => n1372, b => n1373, outb => n5293);
   U4301 : xor2 port map( a => mult_125_G2_ab_6_10_port, b => n1375, outb => 
                           n2923);
   U4302 : xor2 port map( a => mult_125_G2_ab_7_10_port, b => n1377, outb => 
                           n5294);
   U4303 : xor2 port map( a => n4256, b => n4257, outb => n5295);
   U4304 : xor2 port map( a => mult_125_G2_ab_9_10_port, b => n1381, outb => 
                           n5296);
   U4305 : xor2 port map( a => n4260, b => n4258, outb => n5297);
   U4306 : xor2 port map( a => mult_125_G2_ab_11_10_port, b => n1385, outb => 
                           n5298);
   U4307 : xor2 port map( a => n4263, b => n4261, outb => n5299);
   U4308 : xor2 port map( a => mult_125_G2_ab_13_10_port, b => n1389, outb => 
                           n5300);
   U4309 : xor2 port map( a => n4266, b => n4264, outb => n5301);
   U4310 : xor2 port map( a => n5364, b => n1393, outb => n5302);
   U4311 : xor2 port map( a => n1396, b => mult_125_G2_ab_2_9_port, outb => 
                           n2927);
   U4312 : xor2 port map( a => n4269, b => n4267, outb => n5303);
   U4313 : xor2 port map( a => mult_125_G2_ab_4_9_port, b => n1400, outb => 
                           n2929);
   U4314 : xor2 port map( a => mult_125_G2_ab_5_9_port, b => n1402, outb => 
                           n5304);
   U4315 : xor2 port map( a => mult_125_G2_ab_6_9_port, b => n1404, outb => 
                           n2932);
   U4316 : xor2 port map( a => mult_125_G2_ab_7_9_port, b => n1406, outb => 
                           n5305);
   U4317 : xor2 port map( a => n4277, b => n4275, outb => n2935);
   U4318 : xor2 port map( a => n4279, b => n4278, outb => n2938);
   U4319 : xor2 port map( a => mult_125_G2_ab_10_9_port, b => n1412, outb => 
                           n2941);
   U4320 : xor2 port map( a => n4282, b => n4280, outb => n2944);
   U4321 : xor2 port map( a => mult_125_G2_ab_12_9_port, b => n1416, outb => 
                           n2947);
   U4322 : xor2 port map( a => n4285, b => n4283, outb => n2950);
   U4323 : xor2 port map( a => mult_125_G2_ab_14_9_port, b => n1420, outb => 
                           n2953);
   U4324 : xor2 port map( a => n1422, b => n1423, outb => n2955);
   U4325 : xor2 port map( a => n1426, b => mult_125_G2_ab_2_8_port, outb => 
                           n2959);
   U4326 : xor2 port map( a => n4289, b => n4287, outb => n5306);
   U4327 : xor2 port map( a => n4291, b => n1430, outb => n2961);
   U4328 : xor2 port map( a => n4293, b => n4292, outb => n5307);
   U4329 : xor2 port map( a => mult_125_G2_ab_6_8_port, b => n1434, outb => 
                           n2964);
   U4330 : xor2 port map( a => n4296, b => n4294, outb => n5308);
   U4331 : xor2 port map( a => mult_125_G2_ab_8_8_port, b => n1438, outb => 
                           n2967);
   U4332 : xor2 port map( a => mult_125_G2_ab_9_8_port, b => n1440, outb => 
                           n5309);
   U4333 : xor2 port map( a => n4300, b => n4301, outb => n5310);
   U4334 : xor2 port map( a => mult_125_G2_ab_11_8_port, b => n1444, outb => 
                           n5311);
   U4335 : xor2 port map( a => n4304, b => n4302, outb => n5312);
   U4336 : xor2 port map( a => mult_125_G2_ab_13_8_port, b => n1448, outb => 
                           n5313);
   U4337 : xor2 port map( a => n4307, b => n4305, outb => n5314);
   U4338 : xor2 port map( a => n5365, b => n1452, outb => n5315);
   U4339 : xor2 port map( a => n1455, b => mult_125_G2_ab_2_7_port, outb => 
                           n2971);
   U4340 : xor2 port map( a => mult_125_G2_ab_3_7_port, b => n1458, outb => 
                           n5316);
   U4341 : xor2 port map( a => n4311, b => n4310, outb => n2973);
   U4342 : xor2 port map( a => mult_125_G2_ab_5_7_port, b => n1462, outb => 
                           n5317);
   U4343 : xor2 port map( a => n4314, b => n4312, outb => n2976);
   U4344 : xor2 port map( a => mult_125_G2_ab_7_7_port, b => n1466, outb => 
                           n5318);
   U4345 : xor2 port map( a => n4317, b => n4315, outb => n2979);
   U4346 : xor2 port map( a => mult_125_G2_ab_9_7_port, b => n1470, outb => 
                           n5319);
   U4347 : xor2 port map( a => n4320, b => n4318, outb => n2982);
   U4348 : xor2 port map( a => n4322, b => n4321, outb => n2985);
   U4349 : xor2 port map( a => mult_125_G2_ab_12_7_port, b => n1476, outb => 
                           n2988);
   U4350 : xor2 port map( a => n4325, b => n4323, outb => n2991);
   U4351 : xor2 port map( a => mult_125_G2_ab_14_7_port, b => n1480, outb => 
                           n2994);
   U4352 : xor2 port map( a => n1482, b => n1483, outb => n2996);
   U4353 : xor2 port map( a => n1486, b => mult_125_G2_ab_2_6_port, outb => 
                           n3000);
   U4354 : xor2 port map( a => n4329, b => n4327, outb => n5320);
   U4355 : xor2 port map( a => mult_125_G2_ab_4_6_port, b => n1490, outb => 
                           n3002);
   U4356 : xor2 port map( a => n1492, b => n1493, outb => n5321);
   U4357 : xor2 port map( a => mult_125_G2_ab_6_6_port, b => n1495, outb => 
                           n3005);
   U4358 : xor2 port map( a => n4334, b => n4332, outb => n5322);
   U4359 : xor2 port map( a => mult_125_G2_ab_8_6_port, b => n1499, outb => 
                           n3008);
   U4360 : xor2 port map( a => n1501, b => n1502, outb => n5323);
   U4361 : xor2 port map( a => mult_125_G2_ab_10_6_port, b => n1504, outb => 
                           n3011);
   U4362 : xor2 port map( a => mult_125_G2_ab_11_6_port, b => n1506, outb => 
                           n5324);
   U4363 : xor2 port map( a => n4340, b => n4341, outb => n5325);
   U4364 : xor2 port map( a => mult_125_G2_ab_13_6_port, b => n1510, outb => 
                           n5326);
   U4365 : xor2 port map( a => n4344, b => n4342, outb => n5327);
   U4366 : xor2 port map( a => n5366, b => n1514, outb => n5328);
   U4367 : xor2 port map( a => n1517, b => mult_125_G2_ab_2_5_port, outb => 
                           n3015);
   U4368 : xor2 port map( a => mult_125_G2_ab_3_5_port, b => n1520, outb => 
                           n5329);
   U4369 : xor2 port map( a => mult_125_G2_ab_4_5_port, b => n1522, outb => 
                           n3017);
   U4370 : xor2 port map( a => mult_125_G2_ab_5_5_port, b => n1524, outb => 
                           n5330);
   U4371 : xor2 port map( a => n1526, b => n1527, outb => n3020);
   U4372 : xor2 port map( a => mult_125_G2_ab_7_5_port, b => n1529, outb => 
                           n5331);
   U4373 : xor2 port map( a => mult_125_G2_ab_8_5_port, b => n1531, outb => 
                           n3023);
   U4374 : xor2 port map( a => mult_125_G2_ab_9_5_port, b => n1533, outb => 
                           n5332);
   U4375 : xor2 port map( a => n4356, b => n4354, outb => n3026);
   U4376 : xor2 port map( a => mult_125_G2_ab_11_5_port, b => n1537, outb => 
                           n5333);
   U4377 : xor2 port map( a => n4359, b => n4357, outb => n3029);
   U4378 : xor2 port map( a => n4361, b => n1541, outb => n3032);
   U4379 : xor2 port map( a => mult_125_G2_ab_14_5_port, b => n1543, outb => 
                           n3035);
   U4380 : xor2 port map( a => n1545, b => n1546, outb => n3037);
   U4381 : xor2 port map( a => n1549, b => mult_125_G2_ab_2_4_port, outb => 
                           n3041);
   U4382 : xor2 port map( a => n4365, b => n4363, outb => n5334);
   U4383 : xor2 port map( a => mult_125_G2_ab_4_4_port, b => n1553, outb => 
                           n3043);
   U4384 : xor2 port map( a => n1555, b => n1556, outb => n5335);
   U4385 : xor2 port map( a => mult_125_G2_ab_6_4_port, b => n1558, outb => 
                           n3046);
   U4386 : xor2 port map( a => n1560, b => n1561, outb => n5336);
   U4387 : xor2 port map( a => mult_125_G2_ab_8_4_port, b => n1563, outb => 
                           n3049);
   U4388 : xor2 port map( a => mult_125_G2_ab_9_4_port, b => n1565, outb => 
                           n5337);
   U4389 : xor2 port map( a => mult_125_G2_ab_10_4_port, b => n1567, outb => 
                           n3052);
   U4390 : xor2 port map( a => n1569, b => n1570, outb => n5338);
   U4391 : xor2 port map( a => mult_125_G2_ab_12_4_port, b => n1572, outb => 
                           n3055);
   U4392 : xor2 port map( a => mult_125_G2_ab_13_4_port, b => n1574, outb => 
                           n5339);
   U4393 : xor2 port map( a => mult_125_G2_ab_14_4_port, b => n1576, outb => 
                           n5340);
   U4394 : xor2 port map( a => mult_125_G2_ab_15_4_port, b => n1579, outb => 
                           n5341);
   U4395 : xor2 port map( a => n1582, b => mult_125_G2_ab_2_3_port, outb => 
                           n3059);
   U4396 : xor2 port map( a => mult_125_G2_ab_3_3_port, b => n1585, outb => 
                           n5342);
   U4397 : xor2 port map( a => mult_125_G2_ab_4_3_port, b => n1587, outb => 
                           n3061);
   U4398 : xor2 port map( a => mult_125_G2_ab_5_3_port, b => n1589, outb => 
                           n5343);
   U4399 : xor2 port map( a => mult_125_G2_ab_6_3_port, b => n1591, outb => 
                           n3064);
   U4400 : xor2 port map( a => mult_125_G2_ab_7_3_port, b => n1593, outb => 
                           n5344);
   U4401 : xor2 port map( a => mult_125_G2_ab_8_3_port, b => n1595, outb => 
                           n3067);
   U4402 : xor2 port map( a => mult_125_G2_ab_9_3_port, b => n1597, outb => 
                           n5345);
   U4403 : xor2 port map( a => mult_125_G2_ab_10_3_port, b => n1599, outb => 
                           n3070);
   U4404 : xor2 port map( a => mult_125_G2_ab_11_3_port, b => n1601, outb => 
                           n5346);
   U4405 : xor2 port map( a => n4394, b => n4392, outb => n3073);
   U4406 : xor2 port map( a => mult_125_G2_ab_13_3_port, b => n1605, outb => 
                           n5347);
   U4407 : xor2 port map( a => mult_125_G2_ab_14_3_port, b => n1607, outb => 
                           n3076);
   U4408 : xor2 port map( a => mult_125_G2_ab_15_3_port, b => n1609, outb => 
                           n3078);
   U4409 : xor2 port map( a => n1612, b => mult_125_G2_ab_2_2_port, outb => 
                           n3082);
   U4410 : xor2 port map( a => n4400, b => n4398, outb => n5348);
   U4411 : xor2 port map( a => mult_125_G2_ab_4_2_port, b => n1616, outb => 
                           n3084);
   U4412 : xor2 port map( a => mult_125_G2_ab_5_2_port, b => n1618, outb => 
                           n5349);
   U4413 : xor2 port map( a => mult_125_G2_ab_6_2_port, b => n1620, outb => 
                           n3087);
   U4414 : xor2 port map( a => n1622, b => n1623, outb => n5350);
   U4415 : xor2 port map( a => mult_125_G2_ab_8_2_port, b => n1625, outb => 
                           n3090);
   U4416 : xor2 port map( a => mult_125_G2_ab_9_2_port, b => n1627, outb => 
                           n5351);
   U4417 : xor2 port map( a => mult_125_G2_ab_10_2_port, b => n1629, outb => 
                           n3093);
   U4418 : xor2 port map( a => mult_125_G2_ab_11_2_port, b => n1631, outb => 
                           n5352);
   U4419 : xor2 port map( a => mult_125_G2_ab_12_2_port, b => n1633, outb => 
                           n3096);
   U4420 : xor2 port map( a => mult_125_G2_ab_13_2_port, b => n1635, outb => 
                           n5353);
   U4421 : xor2 port map( a => mult_125_G2_ab_14_2_port, b => n1637, outb => 
                           n3099);
   U4422 : xor2 port map( a => n5250, b => n4415, outb => n5354);
   U4423 : xor2 port map( a => n4418, b => mult_125_G2_ab_2_1_port, outb => 
                           n3103);
   U4424 : xor2 port map( a => n4419, b => n4417, outb => n5355);
   U4425 : xor2 port map( a => mult_125_G2_ab_4_1_port, b => n4421, outb => 
                           n3105);
   U4426 : xor2 port map( a => mult_125_G2_ab_5_1_port, b => n1648, outb => 
                           n5367);
   U4427 : xor2 port map( a => n4424, b => n1650, outb => n3108);
   U4428 : xor2 port map( a => n5368, b => n1652, outb => n5357);
   U4429 : xor2 port map( a => mult_125_G2_ab_8_1_port, b => n4425, outb => 
                           n3111);
   U4430 : xor2 port map( a => n5369, b => n1656, outb => n5358);
   U4431 : xor2 port map( a => n4430, b => n1658, outb => n3114);
   U4432 : xor2 port map( a => n5370, b => n1660, outb => n5359);
   U4433 : xor2 port map( a => n4433, b => n1662, outb => n3117);
   U4434 : xor2 port map( a => n5371, b => n1664, outb => n5360);
   U4435 : xor2 port map( a => n4436, b => n4434, outb => n3120);
   U4436 : xor2 port map( a => n5372, b => n1668, outb => n5361);
   U4437 : xor2 port map( a => mult_125_G2_ab_15_0_port, b => n1696, outb => 
                           n5362);
   U4438 : xor2 port map( a => mult_125_G2_ab_11_0_port, b => n1688, outb => 
                           n3122);
   U4439 : xor2 port map( a => mult_125_G2_ab_9_0_port, b => n1684, outb => 
                           n3123);
   U4440 : xor2 port map( a => mult_125_G2_ab_7_0_port, b => n1680, outb => 
                           n3124);
   U4441 : xor2 port map( a => mult_125_G2_ab_5_0_port, b => n1676, outb => 
                           n3125);
   U4442 : xor2 port map( a => mult_125_G2_ab_3_0_port, b => n1672, outb => 
                           n3126);
   U4443 : xor2 port map( a => n344, b => mult_125_G2_ZA, outb => n3127);
   U4444 : xor2 port map( a => mult_125_G2_ab_13_0_port, b => n1692, outb => 
                           n3128);
   U4445 : xor2 port map( a => n5270, b => adder_mem_array_2_32_port, outb => 
                           n3485);
   U4446 : xor2 port map( a => n4808, b => adder_mem_array_2_30_port, outb => 
                           n3487);
   U4447 : xor2 port map( a => n4806, b => adder_mem_array_2_28_port, outb => 
                           n3491);
   U4448 : xor2 port map( a => n4804, b => adder_mem_array_2_26_port, outb => 
                           n3495);
   U4449 : xor2 port map( a => n4802, b => adder_mem_array_2_24_port, outb => 
                           n3499);
   U4450 : xor2 port map( a => n4800, b => adder_mem_array_2_22_port, outb => 
                           n3503);
   U4451 : xor2 port map( a => n4798, b => adder_mem_array_2_20_port, outb => 
                           n3507);
   U4452 : xor2 port map( a => n4796, b => adder_mem_array_2_18_port, outb => 
                           n3511);
   U4453 : xor2 port map( a => n4794, b => adder_mem_array_2_16_port, outb => 
                           n3515);
   U4454 : xor2 port map( a => n4792, b => adder_mem_array_2_14_port, outb => 
                           n3519);
   U4455 : xor2 port map( a => n4790, b => adder_mem_array_2_12_port, outb => 
                           n3523);
   U4456 : xor2 port map( a => n4788, b => adder_mem_array_2_10_port, outb => 
                           n3527);
   U4457 : xor2 port map( a => n4786, b => adder_mem_array_2_8_port, outb => 
                           n3531);
   U4458 : xor2 port map( a => n4784, b => adder_mem_array_2_6_port, outb => 
                           n3535);
   U4459 : xor2 port map( a => n4782, b => adder_mem_array_2_4_port, outb => 
                           n3539);
   U4460 : xor2 port map( a => n4780, b => adder_mem_array_2_2_port, outb => 
                           n3543);
   U4461 : oai22 port map( a => n5374, b => n5375, c => n1698, d => n4464, outb
                           => n5373);
   U4462 : aoi22 port map( a => mult_125_ab_2_15_port, b => 
                           mult_125_ab_3_14_port, c => n5373, d => n5377, outb 
                           => n5376);
   U4463 : oai22 port map( a => n4465, b => n4466, c => n5376, d => n1700, outb
                           => n5378);
   U4464 : aoi22 port map( a => mult_125_ab_4_15_port, b => 
                           mult_125_ab_5_14_port, c => n5378, d => n5380, outb 
                           => n5379);
   U4465 : oai22 port map( a => n4467, b => n4468, c => n5379, d => n1702, outb
                           => n5381);
   U4466 : aoi22 port map( a => mult_125_ab_6_15_port, b => 
                           mult_125_ab_7_14_port, c => n5381, d => n5383, outb 
                           => n5382);
   U4467 : oai22 port map( a => n4469, b => n4470, c => n5382, d => n1704, outb
                           => n5384);
   U4468 : aoi22 port map( a => mult_125_ab_8_15_port, b => 
                           mult_125_ab_9_14_port, c => n5384, d => n5386, outb 
                           => n5385);
   U4469 : oai22 port map( a => n4471, b => n4472, c => n5385, d => n1706, outb
                           => n5387);
   U4470 : aoi22 port map( a => mult_125_ab_10_15_port, b => 
                           mult_125_ab_11_14_port, c => n5387, d => n5389, outb
                           => n5388);
   U4471 : oai22 port map( a => n4473, b => n4474, c => n5388, d => n1708, outb
                           => n5390);
   U4472 : aoi22 port map( a => mult_125_ab_12_15_port, b => 
                           mult_125_ab_13_14_port, c => n5390, d => n5392, outb
                           => n5391);
   U4473 : aoi22 port map( a => mult_125_ab_13_15_port, b => 
                           mult_125_ab_14_14_port, c => n5394, d => n5395, outb
                           => n5393);
   U4474 : aoi22 port map( a => mult_125_ab_14_15_port, b => 
                           mult_125_ab_15_14_port, c => n5396, d => n5397, outb
                           => n277);
   U4475 : inv port map( inb => n4492, outb => n1741);
   U4476 : aoi22 port map( a => n1741, b => mult_125_ab_15_13_port, c => n5398,
                           d => n3171, outb => n279);
   U4477 : aoi22 port map( a => n1770, b => mult_125_ab_15_12_port, c => n5399,
                           d => n3167, outb => n281);
   U4478 : oai22 port map( a => n1801, b => n1800, c => n5401, d => n3212, outb
                           => n5400);
   U4479 : inv port map( inb => n1817, outb => n4542);
   U4480 : aoi22 port map( a => n1831, b => mult_125_ab_15_10_port, c => n5402,
                           d => n3208, outb => n285);
   U4481 : oai22 port map( a => n1861, b => n1860, c => n5404, d => n3253, outb
                           => n5403);
   U4482 : inv port map( inb => n1880, outb => n4586);
   U4483 : aoi22 port map( a => n1890, b => mult_125_ab_15_8_port, c => n5405, 
                           d => n3249, outb => n289);
   U4484 : oai22 port map( a => n1921, b => n1920, c => n5407, d => n3294, outb
                           => n5406);
   U4485 : inv port map( inb => n1946, outb => n4626);
   U4486 : aoi22 port map( a => n1952, b => mult_125_ab_15_6_port, c => n5408, 
                           d => n3290, outb => n293);
   U4487 : oai22 port map( a => n1984, b => n1983, c => n5410, d => n3335, outb
                           => n5409);
   U4488 : aoi22 port map( a => n5411, b => mult_125_ab_15_4_port, c => n2015, 
                           d => n3331, outb => n297);
   U4489 : aoi22 port map( a => n2047, b => mult_125_ab_15_3_port, c => n5412, 
                           d => n3376, outb => n299);
   U4490 : oai22 port map( a => n4700, b => n5413, c => n2076, d => n3372, outb
                           => n302);
   U4491 : aoi22 port map( a => n2106, b => mult_125_ab_15_1_port, c => n5414, 
                           d => n3395, outb => n304);
   U4492 : aoi22 port map( a => n2134, b => mult_125_ab_15_0_port, c => n5415, 
                           d => n5416, outb => n306);
   U4493 : aoi22 port map( a => adder_mem_array_1_1_port, b => n2164, c => 
                           n5417, d => n3447, outb => n3471);
   U4494 : oai22 port map( a => n4777, b => n4778, c => n3471, d => n2165, outb
                           => n3448);
   U4495 : aoi22 port map( a => adder_mem_array_1_3_port, b => 
                           multiplier_sigs_0_3_port, c => n3448, d => n5418, 
                           outb => n3608);
   U4496 : oai22 port map( a => n4810, b => n4811, c => n3608, d => n2201, outb
                           => n3597);
   U4497 : aoi22 port map( a => multiplier_sigs_0_5_port, b => 
                           adder_mem_array_1_5_port, c => n3597, d => n5419, 
                           outb => n3596);
   U4498 : oai22 port map( a => n4812, b => n4813, c => n3596, d => n2203, outb
                           => n3593);
   U4499 : aoi22 port map( a => multiplier_sigs_0_7_port, b => 
                           adder_mem_array_1_7_port, c => n3593, d => n5420, 
                           outb => n3592);
   U4500 : oai22 port map( a => n4814, b => n4815, c => n3592, d => n2205, outb
                           => n3589);
   U4501 : aoi22 port map( a => multiplier_sigs_0_9_port, b => 
                           adder_mem_array_1_9_port, c => n3589, d => n5421, 
                           outb => n3588);
   U4502 : oai22 port map( a => n4816, b => n4817, c => n3588, d => n2207, outb
                           => n3585);
   U4503 : aoi22 port map( a => multiplier_sigs_0_11_port, b => 
                           adder_mem_array_1_11_port, c => n3585, d => n5422, 
                           outb => n3584);
   U4504 : oai22 port map( a => n4818, b => n4819, c => n3584, d => n2209, outb
                           => n3581);
   U4505 : aoi22 port map( a => multiplier_sigs_0_13_port, b => 
                           adder_mem_array_1_13_port, c => n3581, d => n5423, 
                           outb => n3580);
   U4506 : oai22 port map( a => n4820, b => n4821, c => n3580, d => n2211, outb
                           => n3577);
   U4507 : aoi22 port map( a => multiplier_sigs_0_15_port, b => 
                           adder_mem_array_1_15_port, c => n3577, d => n5424, 
                           outb => n3576);
   U4508 : oai22 port map( a => n4822, b => n4823, c => n3576, d => n2213, outb
                           => n3573);
   U4509 : aoi22 port map( a => multiplier_sigs_0_17_port, b => 
                           adder_mem_array_1_17_port, c => n3573, d => n5425, 
                           outb => n3572);
   U4510 : oai22 port map( a => n4824, b => n4825, c => n3572, d => n2215, outb
                           => n3569);
   U4511 : aoi22 port map( a => multiplier_sigs_0_19_port, b => 
                           adder_mem_array_1_19_port, c => n3569, d => n5426, 
                           outb => n3568);
   U4512 : oai22 port map( a => n4826, b => n4827, c => n3568, d => n2217, outb
                           => n3565);
   U4513 : aoi22 port map( a => multiplier_sigs_0_21_port, b => 
                           adder_mem_array_1_21_port, c => n3565, d => n5427, 
                           outb => n3564);
   U4514 : oai22 port map( a => n4828, b => n4829, c => n3564, d => n2219, outb
                           => n3561);
   U4515 : aoi22 port map( a => multiplier_sigs_0_23_port, b => 
                           adder_mem_array_1_23_port, c => n3561, d => n5428, 
                           outb => n3560);
   U4516 : oai22 port map( a => n4830, b => n4831, c => n3560, d => n2221, outb
                           => n3557);
   U4517 : aoi22 port map( a => multiplier_sigs_0_25_port, b => 
                           adder_mem_array_1_25_port, c => n3557, d => n5429, 
                           outb => n3556);
   U4518 : oai22 port map( a => n4832, b => n4833, c => n3556, d => n2223, outb
                           => n3553);
   U4519 : aoi22 port map( a => multiplier_sigs_0_27_port, b => 
                           adder_mem_array_1_27_port, c => n3553, d => n5430, 
                           outb => n3552);
   U4520 : oai22 port map( a => n4834, b => n4835, c => n3552, d => n2225, outb
                           => n3549);
   U4521 : aoi22 port map( a => multiplier_sigs_0_29_port, b => 
                           adder_mem_array_1_29_port, c => n3549, d => n5431, 
                           outb => n3548);
   U4522 : oai22 port map( a => n4836, b => n4837, c => n3548, d => n2227, outb
                           => n2230);
   U4523 : nand2 port map( a => n5432, b => n5433, outb => n2229);
   U4524 : xor2 port map( a => n5373, b => n4894, outb => n3139);
   U4525 : xor2 port map( a => n5434, b => n5376, outb => n3142);
   U4526 : xor2 port map( a => n5378, b => n4895, outb => n3145);
   U4527 : xor2 port map( a => n5435, b => n5379, outb => n3148);
   U4528 : xor2 port map( a => n5381, b => n4896, outb => n3151);
   U4529 : xor2 port map( a => n5436, b => n5382, outb => n3154);
   U4530 : xor2 port map( a => n5384, b => n4897, outb => n3157);
   U4531 : xor2 port map( a => n5437, b => n5385, outb => n3160);
   U4532 : xor2 port map( a => n5387, b => n4898, outb => n3163);
   U4533 : xor2 port map( a => n5438, b => n5388, outb => n3166);
   U4534 : xor2 port map( a => n5390, b => n4899, outb => n3169);
   U4535 : xor2 port map( a => n5439, b => n5394, outb => n3171);
   U4536 : xor2 port map( a => n5393, b => n4900, outb => n280);
   U4537 : xor2 port map( a => n5440, b => n3132, outb => n3177);
   U4538 : xor2 port map( a => n5441, b => n3135, outb => n3183);
   U4539 : xor2 port map( a => n5442, b => n3137, outb => n3186);
   U4540 : xor2 port map( a => n5443, b => n3140, outb => n3189);
   U4541 : xor2 port map( a => n5444, b => n3143, outb => n3192);
   U4542 : xor2 port map( a => n5445, b => n3146, outb => n3195);
   U4543 : xor2 port map( a => n5446, b => n3149, outb => n3198);
   U4544 : xor2 port map( a => n5447, b => n3152, outb => n3201);
   U4545 : xor2 port map( a => n5448, b => n3155, outb => n3204);
   U4546 : xor2 port map( a => n5449, b => n3158, outb => n3207);
   U4547 : xor2 port map( a => n5450, b => n3161, outb => n3210);
   U4548 : xor2 port map( a => n5451, b => n3164, outb => n3212);
   U4549 : xor2 port map( a => n5452, b => n3167, outb => n284);
   U4550 : xor2 port map( a => n5453, b => n3173, outb => n3218);
   U4551 : xor2 port map( a => n5454, b => n3175, outb => n3221);
   U4552 : xor2 port map( a => n5455, b => n3179, outb => n3227);
   U4553 : xor2 port map( a => n5456, b => n3181, outb => n3230);
   U4554 : xor2 port map( a => n5457, b => n3184, outb => n3233);
   U4555 : xor2 port map( a => n5458, b => n3187, outb => n3236);
   U4556 : xor2 port map( a => n5459, b => n3190, outb => n3239);
   U4557 : xor2 port map( a => n5460, b => n3193, outb => n3242);
   U4558 : xor2 port map( a => n5461, b => n3196, outb => n3245);
   U4559 : xor2 port map( a => n5462, b => n3199, outb => n3248);
   U4560 : xor2 port map( a => n5463, b => n3202, outb => n3251);
   U4561 : xor2 port map( a => n5464, b => n3205, outb => n3253);
   U4562 : xor2 port map( a => n5465, b => n3208, outb => n288);
   U4563 : xor2 port map( a => n5466, b => n3214, outb => n3259);
   U4564 : xor2 port map( a => n5467, b => n3216, outb => n3262);
   U4565 : xor2 port map( a => n5468, b => n3219, outb => n3265);
   U4566 : xor2 port map( a => n5469, b => n3223, outb => n3271);
   U4567 : xor2 port map( a => n5470, b => n3225, outb => n3274);
   U4568 : xor2 port map( a => n5471, b => n3228, outb => n3277);
   U4569 : xor2 port map( a => n5472, b => n3231, outb => n3280);
   U4570 : xor2 port map( a => n5473, b => n3234, outb => n3283);
   U4571 : xor2 port map( a => n5474, b => n3237, outb => n3286);
   U4572 : xor2 port map( a => n5475, b => n3240, outb => n3289);
   U4573 : xor2 port map( a => n5476, b => n3243, outb => n3292);
   U4574 : xor2 port map( a => n5477, b => n3246, outb => n3294);
   U4575 : xor2 port map( a => n5478, b => n3249, outb => n292);
   U4576 : xor2 port map( a => n5479, b => n3255, outb => n3300);
   U4577 : xor2 port map( a => n5480, b => n3257, outb => n3303);
   U4578 : xor2 port map( a => n5481, b => n3260, outb => n3306);
   U4579 : xor2 port map( a => n5482, b => n3263, outb => n3309);
   U4580 : xor2 port map( a => n5483, b => n3267, outb => n3315);
   U4581 : xor2 port map( a => n5484, b => n3269, outb => n3318);
   U4582 : xor2 port map( a => n5485, b => n3272, outb => n3321);
   U4583 : xor2 port map( a => n5486, b => n3275, outb => n3324);
   U4584 : xor2 port map( a => n5487, b => n3278, outb => n3327);
   U4585 : xor2 port map( a => n5488, b => n3281, outb => n3330);
   U4586 : xor2 port map( a => n5489, b => n3284, outb => n3333);
   U4587 : xor2 port map( a => n5490, b => n3287, outb => n3335);
   U4588 : xor2 port map( a => n5491, b => n3290, outb => n296);
   U4589 : xor2 port map( a => n5492, b => n3296, outb => n3341);
   U4590 : xor2 port map( a => n5493, b => n3298, outb => n3344);
   U4591 : xor2 port map( a => n5494, b => n3301, outb => n3347);
   U4592 : xor2 port map( a => n5495, b => n3304, outb => n3350);
   U4593 : xor2 port map( a => n5496, b => n3307, outb => n3353);
   U4594 : xor2 port map( a => n5497, b => n3311, outb => n3359);
   U4595 : xor2 port map( a => n5498, b => n3313, outb => n3362);
   U4596 : xor2 port map( a => n5499, b => n3316, outb => n3365);
   U4597 : xor2 port map( a => n5500, b => n3319, outb => n3368);
   U4598 : xor2 port map( a => n5501, b => n3322, outb => n3371);
   U4599 : xor2 port map( a => n5502, b => n3325, outb => n3374);
   U4600 : xor2 port map( a => n5503, b => n3328, outb => n3376);
   U4601 : xor2 port map( a => n5504, b => n3331, outb => n300);
   U4602 : xor2 port map( a => n5505, b => n3337, outb => n3382);
   U4603 : xor2 port map( a => n5506, b => n3339, outb => n3385);
   U4604 : xor2 port map( a => n5507, b => n3342, outb => n3388);
   U4605 : xor2 port map( a => n5508, b => n3345, outb => n3391);
   U4606 : xor2 port map( a => n5509, b => n3348, outb => n3394);
   U4607 : xor2 port map( a => n5510, b => n3351, outb => n3397);
   U4608 : xor2 port map( a => n5511, b => n3355, outb => n3403);
   U4609 : xor2 port map( a => n5512, b => n3357, outb => n3406);
   U4610 : xor2 port map( a => n5513, b => n3360, outb => n3409);
   U4611 : xor2 port map( a => n5514, b => n3363, outb => n3412);
   U4612 : xor2 port map( a => n5515, b => n3366, outb => n3415);
   U4613 : xor2 port map( a => n5516, b => n3369, outb => n3418);
   U4614 : xor2 port map( a => n5517, b => n3372, outb => n305);
   U4615 : xor2 port map( a => n5518, b => n3378, outb => n4728);
   U4616 : xor2 port map( a => n5519, b => n3380, outb => n4732);
   U4617 : xor2 port map( a => n5520, b => n3383, outb => n4736);
   U4618 : xor2 port map( a => n5521, b => n3386, outb => n4740);
   U4619 : xor2 port map( a => n5522, b => n3389, outb => n4744);
   U4620 : xor2 port map( a => n5523, b => n3392, outb => n4748);
   U4621 : inv port map( inb => n3416, outb => n5416);
   U4622 : xor2 port map( a => n5524, b => n3395, outb => n307);
   U4623 : xor2 port map( a => n5525, b => n3416, outb => n311);
   U4624 : xor2 port map( a => n4464, b => mult_125_ab_2_14_port, outb => n3133
                           );
   U4625 : xor2 port map( a => n4465, b => n4466, outb => n5434);
   U4626 : xor2 port map( a => n4467, b => n4468, outb => n5435);
   U4627 : xor2 port map( a => n4469, b => n4470, outb => n5436);
   U4628 : xor2 port map( a => n4471, b => n4472, outb => n5437);
   U4629 : xor2 port map( a => n4473, b => n4474, outb => n5438);
   U4630 : xor2 port map( a => mult_125_ab_13_15_port, b => 
                           mult_125_ab_14_14_port, outb => n5439);
   U4631 : xor2 port map( a => n4475, b => n1713, outb => n3136);
   U4632 : xor2 port map( a => mult_125_ab_3_13_port, b => n1717, outb => n5440
                           );
   U4633 : xor2 port map( a => mult_125_ab_4_13_port, b => n1719, outb => n3138
                           );
   U4634 : xor2 port map( a => mult_125_ab_5_13_port, b => n1721, outb => n3141
                           );
   U4635 : xor2 port map( a => mult_125_ab_6_13_port, b => n1723, outb => n3144
                           );
   U4636 : xor2 port map( a => n4482, b => n4480, outb => n3147);
   U4637 : xor2 port map( a => mult_125_ab_8_13_port, b => n1727, outb => n3150
                           );
   U4638 : xor2 port map( a => n4485, b => n4483, outb => n3153);
   U4639 : xor2 port map( a => mult_125_ab_10_13_port, b => n1731, outb => 
                           n3156);
   U4640 : xor2 port map( a => n4488, b => n4486, outb => n3159);
   U4641 : xor2 port map( a => mult_125_ab_12_13_port, b => n1735, outb => 
                           n3162);
   U4642 : xor2 port map( a => n4491, b => n4489, outb => n3165);
   U4643 : xor2 port map( a => mult_125_ab_14_13_port, b => n1739, outb => 
                           n3168);
   U4644 : xor2 port map( a => mult_125_ab_15_13_port, b => n4492, outb => 
                           n3170);
   U4645 : xor2 port map( a => n1744, b => mult_125_ab_2_12_port, outb => n3174
                           );
   U4646 : xor2 port map( a => n4496, b => n4494, outb => n5441);
   U4647 : xor2 port map( a => mult_125_ab_4_12_port, b => n1748, outb => n3176
                           );
   U4648 : xor2 port map( a => mult_125_ab_5_12_port, b => n4497, outb => n5442
                           );
   U4649 : xor2 port map( a => n4501, b => n4499, outb => n5443);
   U4650 : xor2 port map( a => mult_125_ab_7_12_port, b => n1754, outb => n5444
                           );
   U4651 : xor2 port map( a => n4504, b => n4502, outb => n5445);
   U4652 : xor2 port map( a => mult_125_ab_9_12_port, b => n1758, outb => n5446
                           );
   U4653 : xor2 port map( a => n4507, b => n4505, outb => n5447);
   U4654 : xor2 port map( a => mult_125_ab_11_12_port, b => n1762, outb => 
                           n5448);
   U4655 : xor2 port map( a => n4510, b => n4508, outb => n5449);
   U4656 : xor2 port map( a => mult_125_ab_13_12_port, b => n1766, outb => 
                           n5450);
   U4657 : xor2 port map( a => n4513, b => n4511, outb => n5451);
   U4658 : xor2 port map( a => n5526, b => n1770, outb => n5452);
   U4659 : xor2 port map( a => n1773, b => mult_125_ab_2_11_port, outb => n3180
                           );
   U4660 : xor2 port map( a => mult_125_ab_3_11_port, b => n1776, outb => n5453
                           );
   U4661 : xor2 port map( a => n4517, b => n4516, outb => n3182);
   U4662 : xor2 port map( a => mult_125_ab_5_11_port, b => n1780, outb => n5454
                           );
   U4663 : xor2 port map( a => mult_125_ab_6_11_port, b => n1782, outb => n3185
                           );
   U4664 : xor2 port map( a => n4522, b => n4521, outb => n3188);
   U4665 : xor2 port map( a => mult_125_ab_8_11_port, b => n1786, outb => n3191
                           );
   U4666 : xor2 port map( a => n4525, b => n4523, outb => n3194);
   U4667 : xor2 port map( a => mult_125_ab_10_11_port, b => n1790, outb => 
                           n3197);
   U4668 : xor2 port map( a => n4528, b => n4526, outb => n3200);
   U4669 : xor2 port map( a => mult_125_ab_12_11_port, b => n1794, outb => 
                           n3203);
   U4670 : xor2 port map( a => n4531, b => n4529, outb => n3206);
   U4671 : xor2 port map( a => mult_125_ab_14_11_port, b => n1798, outb => 
                           n3209);
   U4672 : xor2 port map( a => n1800, b => n1801, outb => n3211);
   U4673 : xor2 port map( a => n1804, b => mult_125_ab_2_10_port, outb => n3215
                           );
   U4674 : xor2 port map( a => n4535, b => n4533, outb => n5455);
   U4675 : xor2 port map( a => mult_125_ab_4_10_port, b => n1808, outb => n3217
                           );
   U4676 : xor2 port map( a => n1810, b => n1811, outb => n5456);
   U4677 : xor2 port map( a => mult_125_ab_6_10_port, b => n1813, outb => n3220
                           );
   U4678 : xor2 port map( a => mult_125_ab_7_10_port, b => n1815, outb => n5457
                           );
   U4679 : xor2 port map( a => n4541, b => n4542, outb => n5458);
   U4680 : xor2 port map( a => mult_125_ab_9_10_port, b => n1819, outb => n5459
                           );
   U4681 : xor2 port map( a => n4545, b => n4543, outb => n5460);
   U4682 : xor2 port map( a => mult_125_ab_11_10_port, b => n1823, outb => 
                           n5461);
   U4683 : xor2 port map( a => n4548, b => n4546, outb => n5462);
   U4684 : xor2 port map( a => mult_125_ab_13_10_port, b => n1827, outb => 
                           n5463);
   U4685 : xor2 port map( a => n4551, b => n4549, outb => n5464);
   U4686 : xor2 port map( a => n5527, b => n1831, outb => n5465);
   U4687 : xor2 port map( a => n1834, b => mult_125_ab_2_9_port, outb => n3224)
                           ;
   U4688 : xor2 port map( a => n4554, b => n4552, outb => n5466);
   U4689 : xor2 port map( a => mult_125_ab_4_9_port, b => n1838, outb => n3226)
                           ;
   U4690 : xor2 port map( a => mult_125_ab_5_9_port, b => n1840, outb => n5467)
                           ;
   U4691 : xor2 port map( a => mult_125_ab_6_9_port, b => n1842, outb => n3229)
                           ;
   U4692 : xor2 port map( a => mult_125_ab_7_9_port, b => n1844, outb => n5468)
                           ;
   U4693 : xor2 port map( a => n4562, b => n4560, outb => n3232);
   U4694 : xor2 port map( a => n4564, b => n4563, outb => n3235);
   U4695 : xor2 port map( a => mult_125_ab_10_9_port, b => n1850, outb => n3238
                           );
   U4696 : xor2 port map( a => n4567, b => n4565, outb => n3241);
   U4697 : xor2 port map( a => mult_125_ab_12_9_port, b => n1854, outb => n3244
                           );
   U4698 : xor2 port map( a => n4570, b => n4568, outb => n3247);
   U4699 : xor2 port map( a => mult_125_ab_14_9_port, b => n1858, outb => n3250
                           );
   U4700 : xor2 port map( a => n1860, b => n1861, outb => n3252);
   U4701 : xor2 port map( a => n1864, b => mult_125_ab_2_8_port, outb => n3256)
                           ;
   U4702 : xor2 port map( a => n4574, b => n4572, outb => n5469);
   U4703 : xor2 port map( a => n4576, b => n1868, outb => n3258);
   U4704 : xor2 port map( a => n4578, b => n4577, outb => n5470);
   U4705 : xor2 port map( a => mult_125_ab_6_8_port, b => n1872, outb => n3261)
                           ;
   U4706 : xor2 port map( a => n4581, b => n4579, outb => n5471);
   U4707 : xor2 port map( a => mult_125_ab_8_8_port, b => n1876, outb => n3264)
                           ;
   U4708 : xor2 port map( a => mult_125_ab_9_8_port, b => n1878, outb => n5472)
                           ;
   U4709 : xor2 port map( a => n4585, b => n4586, outb => n5473);
   U4710 : xor2 port map( a => mult_125_ab_11_8_port, b => n1882, outb => n5474
                           );
   U4711 : xor2 port map( a => n4589, b => n4587, outb => n5475);
   U4712 : xor2 port map( a => mult_125_ab_13_8_port, b => n1886, outb => n5476
                           );
   U4713 : xor2 port map( a => n4592, b => n4590, outb => n5477);
   U4714 : xor2 port map( a => n5528, b => n1890, outb => n5478);
   U4715 : xor2 port map( a => n1893, b => mult_125_ab_2_7_port, outb => n3268)
                           ;
   U4716 : xor2 port map( a => mult_125_ab_3_7_port, b => n1896, outb => n5479)
                           ;
   U4717 : xor2 port map( a => n4596, b => n4595, outb => n3270);
   U4718 : xor2 port map( a => mult_125_ab_5_7_port, b => n1900, outb => n5480)
                           ;
   U4719 : xor2 port map( a => n4599, b => n4597, outb => n3273);
   U4720 : xor2 port map( a => mult_125_ab_7_7_port, b => n1904, outb => n5481)
                           ;
   U4721 : xor2 port map( a => n4602, b => n4600, outb => n3276);
   U4722 : xor2 port map( a => mult_125_ab_9_7_port, b => n1908, outb => n5482)
                           ;
   U4723 : xor2 port map( a => n4605, b => n4603, outb => n3279);
   U4724 : xor2 port map( a => n4607, b => n4606, outb => n3282);
   U4725 : xor2 port map( a => mult_125_ab_12_7_port, b => n1914, outb => n3285
                           );
   U4726 : xor2 port map( a => n4610, b => n4608, outb => n3288);
   U4727 : xor2 port map( a => mult_125_ab_14_7_port, b => n1918, outb => n3291
                           );
   U4728 : xor2 port map( a => n1920, b => n1921, outb => n3293);
   U4729 : xor2 port map( a => n1924, b => mult_125_ab_2_6_port, outb => n3297)
                           ;
   U4730 : xor2 port map( a => n4614, b => n4612, outb => n5483);
   U4731 : xor2 port map( a => mult_125_ab_4_6_port, b => n1928, outb => n3299)
                           ;
   U4732 : xor2 port map( a => n1930, b => n1931, outb => n5484);
   U4733 : xor2 port map( a => mult_125_ab_6_6_port, b => n1933, outb => n3302)
                           ;
   U4734 : xor2 port map( a => n4619, b => n4617, outb => n5485);
   U4735 : xor2 port map( a => mult_125_ab_8_6_port, b => n1937, outb => n3305)
                           ;
   U4736 : xor2 port map( a => n1939, b => n1940, outb => n5486);
   U4737 : xor2 port map( a => mult_125_ab_10_6_port, b => n1942, outb => n3308
                           );
   U4738 : xor2 port map( a => mult_125_ab_11_6_port, b => n1944, outb => n5487
                           );
   U4739 : xor2 port map( a => n4625, b => n4626, outb => n5488);
   U4740 : xor2 port map( a => mult_125_ab_13_6_port, b => n1948, outb => n5489
                           );
   U4741 : xor2 port map( a => n4629, b => n4627, outb => n5490);
   U4742 : xor2 port map( a => n5529, b => n1952, outb => n5491);
   U4743 : xor2 port map( a => n1955, b => mult_125_ab_2_5_port, outb => n3312)
                           ;
   U4744 : xor2 port map( a => mult_125_ab_3_5_port, b => n1958, outb => n5492)
                           ;
   U4745 : xor2 port map( a => mult_125_ab_4_5_port, b => n1960, outb => n3314)
                           ;
   U4746 : xor2 port map( a => mult_125_ab_5_5_port, b => n1962, outb => n5493)
                           ;
   U4747 : xor2 port map( a => n1964, b => n1965, outb => n3317);
   U4748 : xor2 port map( a => mult_125_ab_7_5_port, b => n1967, outb => n5494)
                           ;
   U4749 : xor2 port map( a => mult_125_ab_8_5_port, b => n1969, outb => n3320)
                           ;
   U4750 : xor2 port map( a => mult_125_ab_9_5_port, b => n1971, outb => n5495)
                           ;
   U4751 : xor2 port map( a => n4641, b => n4639, outb => n3323);
   U4752 : xor2 port map( a => mult_125_ab_11_5_port, b => n1975, outb => n5496
                           );
   U4753 : xor2 port map( a => n4644, b => n4642, outb => n3326);
   U4754 : xor2 port map( a => n4646, b => n1979, outb => n3329);
   U4755 : xor2 port map( a => mult_125_ab_14_5_port, b => n1981, outb => n3332
                           );
   U4756 : xor2 port map( a => n1983, b => n1984, outb => n3334);
   U4757 : xor2 port map( a => n1987, b => mult_125_ab_2_4_port, outb => n3338)
                           ;
   U4758 : xor2 port map( a => n4650, b => n4648, outb => n5497);
   U4759 : xor2 port map( a => mult_125_ab_4_4_port, b => n1991, outb => n3340)
                           ;
   U4760 : xor2 port map( a => n1993, b => n1994, outb => n5498);
   U4761 : xor2 port map( a => mult_125_ab_6_4_port, b => n1996, outb => n3343)
                           ;
   U4762 : xor2 port map( a => n1998, b => n1999, outb => n5499);
   U4763 : xor2 port map( a => mult_125_ab_8_4_port, b => n2001, outb => n3346)
                           ;
   U4764 : xor2 port map( a => mult_125_ab_9_4_port, b => n2003, outb => n5500)
                           ;
   U4765 : xor2 port map( a => mult_125_ab_10_4_port, b => n2005, outb => n3349
                           );
   U4766 : xor2 port map( a => n2007, b => n2008, outb => n5501);
   U4767 : xor2 port map( a => mult_125_ab_12_4_port, b => n2010, outb => n3352
                           );
   U4768 : xor2 port map( a => mult_125_ab_13_4_port, b => n2012, outb => n5502
                           );
   U4769 : xor2 port map( a => mult_125_ab_14_4_port, b => n2014, outb => n5503
                           );
   U4770 : xor2 port map( a => mult_125_ab_15_4_port, b => n2017, outb => n5504
                           );
   U4771 : xor2 port map( a => n2020, b => mult_125_ab_2_3_port, outb => n3356)
                           ;
   U4772 : xor2 port map( a => mult_125_ab_3_3_port, b => n2023, outb => n5505)
                           ;
   U4773 : xor2 port map( a => mult_125_ab_4_3_port, b => n2025, outb => n3358)
                           ;
   U4774 : xor2 port map( a => mult_125_ab_5_3_port, b => n2027, outb => n5506)
                           ;
   U4775 : xor2 port map( a => mult_125_ab_6_3_port, b => n2029, outb => n3361)
                           ;
   U4776 : xor2 port map( a => mult_125_ab_7_3_port, b => n2031, outb => n5507)
                           ;
   U4777 : xor2 port map( a => mult_125_ab_8_3_port, b => n2033, outb => n3364)
                           ;
   U4778 : xor2 port map( a => mult_125_ab_9_3_port, b => n2035, outb => n5508)
                           ;
   U4779 : xor2 port map( a => mult_125_ab_10_3_port, b => n2037, outb => n3367
                           );
   U4780 : xor2 port map( a => mult_125_ab_11_3_port, b => n2039, outb => n5509
                           );
   U4781 : xor2 port map( a => n4679, b => n4677, outb => n3370);
   U4782 : xor2 port map( a => mult_125_ab_13_3_port, b => n2043, outb => n5510
                           );
   U4783 : xor2 port map( a => mult_125_ab_14_3_port, b => n2045, outb => n3373
                           );
   U4784 : xor2 port map( a => mult_125_ab_15_3_port, b => n2047, outb => n3375
                           );
   U4785 : xor2 port map( a => n2050, b => mult_125_ab_2_2_port, outb => n3379)
                           ;
   U4786 : xor2 port map( a => n4685, b => n4683, outb => n5511);
   U4787 : xor2 port map( a => mult_125_ab_4_2_port, b => n2054, outb => n3381)
                           ;
   U4788 : xor2 port map( a => mult_125_ab_5_2_port, b => n2056, outb => n5512)
                           ;
   U4789 : xor2 port map( a => mult_125_ab_6_2_port, b => n2058, outb => n3384)
                           ;
   U4790 : xor2 port map( a => n2060, b => n2061, outb => n5513);
   U4791 : xor2 port map( a => mult_125_ab_8_2_port, b => n2063, outb => n3387)
                           ;
   U4792 : xor2 port map( a => mult_125_ab_9_2_port, b => n2065, outb => n5514)
                           ;
   U4793 : xor2 port map( a => mult_125_ab_10_2_port, b => n2067, outb => n3390
                           );
   U4794 : xor2 port map( a => mult_125_ab_11_2_port, b => n2069, outb => n5515
                           );
   U4795 : xor2 port map( a => mult_125_ab_12_2_port, b => n2071, outb => n3393
                           );
   U4796 : xor2 port map( a => mult_125_ab_13_2_port, b => n2073, outb => n5516
                           );
   U4797 : xor2 port map( a => mult_125_ab_14_2_port, b => n2075, outb => n3396
                           );
   U4798 : xor2 port map( a => n5413, b => n4700, outb => n5517);
   U4799 : xor2 port map( a => n4703, b => mult_125_ab_2_1_port, outb => n3400)
                           ;
   U4800 : xor2 port map( a => n4704, b => n4702, outb => n5518);
   U4801 : xor2 port map( a => mult_125_ab_4_1_port, b => n4706, outb => n3402)
                           ;
   U4802 : xor2 port map( a => mult_125_ab_5_1_port, b => n2086, outb => n5530)
                           ;
   U4803 : xor2 port map( a => n4709, b => n2088, outb => n3405);
   U4804 : xor2 port map( a => n5531, b => n2090, outb => n5520);
   U4805 : xor2 port map( a => mult_125_ab_8_1_port, b => n4710, outb => n3408)
                           ;
   U4806 : xor2 port map( a => n5532, b => n2094, outb => n5521);
   U4807 : xor2 port map( a => n4715, b => n2096, outb => n3411);
   U4808 : xor2 port map( a => n5533, b => n2098, outb => n5522);
   U4809 : xor2 port map( a => n4718, b => n2100, outb => n3414);
   U4810 : xor2 port map( a => n5534, b => n2102, outb => n5523);
   U4811 : xor2 port map( a => n4721, b => n4719, outb => n3417);
   U4812 : xor2 port map( a => n5535, b => n2106, outb => n5524);
   U4813 : xor2 port map( a => mult_125_ab_15_0_port, b => n2134, outb => n5525
                           );
   U4814 : xor2 port map( a => mult_125_ab_11_0_port, b => n2126, outb => n3419
                           );
   U4815 : xor2 port map( a => mult_125_ab_9_0_port, b => n2122, outb => n3420)
                           ;
   U4816 : xor2 port map( a => mult_125_ab_7_0_port, b => n2118, outb => n3421)
                           ;
   U4817 : xor2 port map( a => mult_125_ab_5_0_port, b => n2114, outb => n3422)
                           ;
   U4818 : xor2 port map( a => mult_125_ab_3_0_port, b => n2110, outb => n3423)
                           ;
   U4819 : xor2 port map( a => n308, b => mult_125_ZA, outb => n3424);
   U4820 : xor2 port map( a => mult_125_ab_13_0_port, b => n2130, outb => n3425
                           );
   U4821 : xor2 port map( a => n4777, b => adder_mem_array_1_2_port, outb => 
                           n3470);
   U4822 : xor2 port map( a => n5433, b => adder_mem_array_1_32_port, outb => 
                           n3545);
   U4823 : xor2 port map( a => n4836, b => adder_mem_array_1_30_port, outb => 
                           n3547);
   U4824 : xor2 port map( a => n4834, b => adder_mem_array_1_28_port, outb => 
                           n3551);
   U4825 : xor2 port map( a => n4832, b => adder_mem_array_1_26_port, outb => 
                           n3555);
   U4826 : xor2 port map( a => n4830, b => adder_mem_array_1_24_port, outb => 
                           n3559);
   U4827 : xor2 port map( a => n4828, b => adder_mem_array_1_22_port, outb => 
                           n3563);
   U4828 : xor2 port map( a => n4826, b => adder_mem_array_1_20_port, outb => 
                           n3567);
   U4829 : xor2 port map( a => n4824, b => adder_mem_array_1_18_port, outb => 
                           n3571);
   U4830 : xor2 port map( a => n4822, b => adder_mem_array_1_16_port, outb => 
                           n3575);
   U4831 : xor2 port map( a => n4820, b => adder_mem_array_1_14_port, outb => 
                           n3579);
   U4832 : xor2 port map( a => n4818, b => adder_mem_array_1_12_port, outb => 
                           n3583);
   U4833 : xor2 port map( a => n4816, b => adder_mem_array_1_10_port, outb => 
                           n3587);
   U4834 : xor2 port map( a => n4814, b => adder_mem_array_1_8_port, outb => 
                           n3591);
   U4835 : xor2 port map( a => n4812, b => adder_mem_array_1_6_port, outb => 
                           n3595);
   U4836 : xor2 port map( a => n4810, b => adder_mem_array_1_4_port, outb => 
                           n3607);
   U4837 : inv port map( inb => n385, outb => n4905);
   U4838 : inv port map( inb => n387, outb => n4908);
   U4839 : inv port map( inb => n389, outb => n4911);
   U4840 : inv port map( inb => n391, outb => n4914);
   U4841 : inv port map( inb => n393, outb => n4917);
   U4842 : inv port map( inb => n395, outb => n4920);
   U4843 : inv port map( inb => n397, outb => n4925);
   U4844 : inv port map( inb => n430, outb => n3640);
   U4845 : inv port map( inb => n459, outb => n3659);
   U4846 : inv port map( inb => n490, outb => n3679);
   U4847 : inv port map( inb => n520, outb => n3698);
   U4848 : inv port map( inb => n550, outb => n3718);
   U4849 : inv port map( inb => n579, outb => n3738);
   U4850 : inv port map( inb => n610, outb => n3758);
   U4851 : inv port map( inb => n641, outb => n3775);
   U4852 : inv port map( inb => n673, outb => n3794);
   U4853 : inv port map( inb => n706, outb => n3809);
   U4854 : inv port map( inb => n736, outb => n3829);
   U4855 : inv port map( inb => n766, outb => n3848);
   U4856 : inv port map( inb => n3867, outb => n794);
   U4857 : inv port map( inb => n3868, outb => n796);
   U4858 : inv port map( inb => n819, outb => n4943);
   U4859 : inv port map( inb => n823, outb => n5051);
   U4860 : inv port map( inb => n825, outb => n5054);
   U4861 : inv port map( inb => n827, outb => n5057);
   U4862 : inv port map( inb => n829, outb => n5060);
   U4863 : inv port map( inb => n831, outb => n5063);
   U4864 : inv port map( inb => n833, outb => n5066);
   U4865 : inv port map( inb => n835, outb => n5071);
   U4866 : inv port map( inb => n868, outb => n3925);
   U4867 : inv port map( inb => n897, outb => n3944);
   U4868 : inv port map( inb => n928, outb => n3964);
   U4869 : inv port map( inb => n958, outb => n3983);
   U4870 : inv port map( inb => n988, outb => n4003);
   U4871 : inv port map( inb => n1017, outb => n4023);
   U4872 : inv port map( inb => n1048, outb => n4043);
   U4873 : inv port map( inb => n1079, outb => n4060);
   U4874 : inv port map( inb => n1111, outb => n4079);
   U4875 : inv port map( inb => n1144, outb => n4094);
   U4876 : inv port map( inb => n1174, outb => n4114);
   U4877 : inv port map( inb => n1204, outb => n4133);
   U4878 : inv port map( inb => n4152, outb => n1232);
   U4879 : inv port map( inb => n4153, outb => n1234);
   U4880 : inv port map( inb => n1257, outb => n5089);
   U4881 : inv port map( inb => n1261, outb => n5214);
   U4882 : inv port map( inb => n1263, outb => n5217);
   U4883 : inv port map( inb => n1265, outb => n5220);
   U4884 : inv port map( inb => n1267, outb => n5223);
   U4885 : inv port map( inb => n1269, outb => n5226);
   U4886 : inv port map( inb => n1271, outb => n5229);
   U4887 : inv port map( inb => n1273, outb => n5234);
   U4888 : inv port map( inb => n1306, outb => n4210);
   U4889 : inv port map( inb => n1335, outb => n4229);
   U4890 : inv port map( inb => n1366, outb => n4249);
   U4891 : inv port map( inb => n1396, outb => n4268);
   U4892 : inv port map( inb => n1426, outb => n4288);
   U4893 : inv port map( inb => n1455, outb => n4308);
   U4894 : inv port map( inb => n1486, outb => n4328);
   U4895 : inv port map( inb => n1517, outb => n4345);
   U4896 : inv port map( inb => n1549, outb => n4364);
   U4897 : inv port map( inb => n1582, outb => n4379);
   U4898 : inv port map( inb => n1612, outb => n4399);
   U4899 : inv port map( inb => n1642, outb => n4418);
   U4900 : inv port map( inb => n4437, outb => n1670);
   U4901 : inv port map( inb => n4438, outb => n1672);
   U4902 : inv port map( inb => n1695, outb => n5252);
   U4903 : inv port map( inb => n1699, outb => n5377);
   U4904 : inv port map( inb => n1701, outb => n5380);
   U4905 : inv port map( inb => n1703, outb => n5383);
   U4906 : inv port map( inb => n1705, outb => n5386);
   U4907 : inv port map( inb => n1707, outb => n5389);
   U4908 : inv port map( inb => n1709, outb => n5392);
   U4909 : inv port map( inb => n1711, outb => n5397);
   U4910 : inv port map( inb => n1744, outb => n4495);
   U4911 : inv port map( inb => n1773, outb => n4514);
   U4912 : inv port map( inb => n1804, outb => n4534);
   U4913 : inv port map( inb => n1834, outb => n4553);
   U4914 : inv port map( inb => n1864, outb => n4573);
   U4915 : inv port map( inb => n1893, outb => n4593);
   U4916 : inv port map( inb => n1924, outb => n4613);
   U4917 : inv port map( inb => n1955, outb => n4630);
   U4918 : inv port map( inb => n1987, outb => n4649);
   U4919 : inv port map( inb => n2020, outb => n4664);
   U4920 : inv port map( inb => n2050, outb => n4684);
   U4921 : inv port map( inb => n2080, outb => n4703);
   U4922 : inv port map( inb => n4722, outb => n2108);
   U4923 : inv port map( inb => n4723, outb => n2110);
   U4924 : inv port map( inb => n2133, outb => n5415);
   U4925 : inv port map( inb => n4749, outb => n2137);
   U4926 : inv port map( inb => n2139, outb => n5092);
   U4927 : inv port map( inb => n2141, outb => n5093);
   U4928 : inv port map( inb => n2143, outb => n5094);
   U4929 : inv port map( inb => n2145, outb => n5095);
   U4930 : inv port map( inb => n2147, outb => n5096);
   U4931 : inv port map( inb => n2149, outb => n5097);
   U4932 : inv port map( inb => n2151, outb => n5098);
   U4933 : inv port map( inb => n2153, outb => n5099);
   U4934 : inv port map( inb => n2155, outb => n5100);
   U4935 : inv port map( inb => n2157, outb => n5101);
   U4936 : inv port map( inb => n2159, outb => n5102);
   U4937 : inv port map( inb => n2161, outb => n5103);
   U4938 : inv port map( inb => n4776, outb => n2164);
   U4939 : inv port map( inb => n4779, outb => n2167);
   U4940 : inv port map( inb => n2169, outb => n5255);
   U4941 : inv port map( inb => n2171, outb => n5256);
   U4942 : inv port map( inb => n2173, outb => n5257);
   U4943 : inv port map( inb => n2175, outb => n5258);
   U4944 : inv port map( inb => n2177, outb => n5259);
   U4945 : inv port map( inb => n2179, outb => n5260);
   U4946 : inv port map( inb => n2181, outb => n5261);
   U4947 : inv port map( inb => n2183, outb => n5262);
   U4948 : inv port map( inb => n2185, outb => n5263);
   U4949 : inv port map( inb => n2187, outb => n5264);
   U4950 : inv port map( inb => n2189, outb => n5265);
   U4951 : inv port map( inb => n2191, outb => n5266);
   U4952 : inv port map( inb => n2193, outb => n5267);
   U4953 : inv port map( inb => n2195, outb => n5268);
   U4954 : inv port map( inb => n2200, outb => n5418);
   U4955 : inv port map( inb => n2202, outb => n5419);
   U4956 : inv port map( inb => n2204, outb => n5420);
   U4957 : inv port map( inb => n2206, outb => n5421);
   U4958 : inv port map( inb => n2208, outb => n5422);
   U4959 : inv port map( inb => n2210, outb => n5423);
   U4960 : inv port map( inb => n2212, outb => n5424);
   U4961 : inv port map( inb => n2214, outb => n5425);
   U4962 : inv port map( inb => n2216, outb => n5426);
   U4963 : inv port map( inb => n2218, outb => n5427);
   U4964 : inv port map( inb => n2220, outb => n5428);
   U4965 : inv port map( inb => n2222, outb => n5429);
   U4966 : inv port map( inb => n2224, outb => n5430);
   U4967 : inv port map( inb => n2226, outb => n5431);
   U4968 : inv port map( inb => n2231, outb => n5104);
   U4969 : inv port map( inb => n2233, outb => n5105);
   U4970 : inv port map( inb => mult_125_G4_ab_1_15_port, outb => n4902);
   U4971 : inv port map( inb => mult_125_G4_ab_2_14_port, outb => n4903);
   U4972 : inv port map( inb => n408, outb => n3626);
   U4973 : inv port map( inb => n412, outb => n3629);
   U4974 : inv port map( inb => n416, outb => n3632);
   U4975 : inv port map( inb => n420, outb => n3635);
   U4976 : inv port map( inb => n424, outb => n3638);
   U4977 : inv port map( inb => mult_125_G4_ab_3_12_port, outb => n3641);
   U4978 : inv port map( inb => n439, outb => n3648);
   U4979 : inv port map( inb => n443, outb => n3651);
   U4980 : inv port map( inb => n447, outb => n3654);
   U4981 : inv port map( inb => n451, outb => n3657);
   U4982 : inv port map( inb => mult_125_G4_ab_3_11_port, outb => n461);
   U4983 : inv port map( inb => n471, outb => n3669);
   U4984 : inv port map( inb => n475, outb => n3672);
   U4985 : inv port map( inb => n479, outb => n3675);
   U4986 : inv port map( inb => n483, outb => n3677);
   U4987 : inv port map( inb => mult_125_G4_ab_3_10_port, outb => n3680);
   U4988 : inv port map( inb => n504, outb => n3689);
   U4989 : inv port map( inb => n508, outb => n3692);
   U4990 : inv port map( inb => n512, outb => n3695);
   U4991 : inv port map( inb => mult_125_G4_ab_3_9_port, outb => n3699);
   U4992 : inv port map( inb => n535, outb => n3711);
   U4993 : inv port map( inb => n539, outb => n3714);
   U4994 : inv port map( inb => n543, outb => n3716);
   U4995 : inv port map( inb => mult_125_G4_ab_3_8_port, outb => n3719);
   U4996 : inv port map( inb => n567, outb => n3733);
   U4997 : inv port map( inb => n571, outb => n3736);
   U4998 : inv port map( inb => mult_125_G4_ab_3_7_port, outb => n581);
   U4999 : inv port map( inb => n599, outb => n3754);
   U5000 : inv port map( inb => n603, outb => n3756);
   U5001 : inv port map( inb => mult_125_G4_ab_3_6_port, outb => n3759);
   U5002 : inv port map( inb => n633, outb => n3773);
   U5003 : inv port map( inb => mult_125_G4_ab_3_5_port, outb => n643);
   U5004 : inv port map( inb => n666, outb => n3792);
   U5005 : inv port map( inb => mult_125_G4_ab_3_4_port, outb => n3795);
   U5006 : inv port map( inb => mult_125_G4_ab_3_3_port, outb => n708);
   U5007 : inv port map( inb => mult_125_G4_ab_3_2_port, outb => n3830);
   U5008 : inv port map( inb => mult_125_G4_ab_3_1_port, outb => n3849);
   U5009 : inv port map( inb => n770, outb => n3851);
   U5010 : inv port map( inb => n799, outb => n3875);
   U5011 : inv port map( inb => n803, outb => n3879);
   U5012 : inv port map( inb => n807, outb => n3883);
   U5013 : inv port map( inb => n811, outb => n3887);
   U5014 : inv port map( inb => n815, outb => n3891);
   U5015 : inv port map( inb => mult_125_G3_ab_1_15_port, outb => n5048);
   U5016 : inv port map( inb => mult_125_G3_ab_2_14_port, outb => n5049);
   U5017 : inv port map( inb => n846, outb => n3911);
   U5018 : inv port map( inb => n850, outb => n3914);
   U5019 : inv port map( inb => n854, outb => n3917);
   U5020 : inv port map( inb => n858, outb => n3920);
   U5021 : inv port map( inb => n862, outb => n3923);
   U5022 : inv port map( inb => mult_125_G3_ab_3_12_port, outb => n3926);
   U5023 : inv port map( inb => n877, outb => n3933);
   U5024 : inv port map( inb => n881, outb => n3936);
   U5025 : inv port map( inb => n885, outb => n3939);
   U5026 : inv port map( inb => n889, outb => n3942);
   U5027 : inv port map( inb => mult_125_G3_ab_3_11_port, outb => n899);
   U5028 : inv port map( inb => n909, outb => n3954);
   U5029 : inv port map( inb => n913, outb => n3957);
   U5030 : inv port map( inb => n917, outb => n3960);
   U5031 : inv port map( inb => n921, outb => n3962);
   U5032 : inv port map( inb => mult_125_G3_ab_3_10_port, outb => n3965);
   U5033 : inv port map( inb => n942, outb => n3974);
   U5034 : inv port map( inb => n946, outb => n3977);
   U5035 : inv port map( inb => n950, outb => n3980);
   U5036 : inv port map( inb => mult_125_G3_ab_3_9_port, outb => n3984);
   U5037 : inv port map( inb => n973, outb => n3996);
   U5038 : inv port map( inb => n977, outb => n3999);
   U5039 : inv port map( inb => n981, outb => n4001);
   U5040 : inv port map( inb => mult_125_G3_ab_3_8_port, outb => n4004);
   U5041 : inv port map( inb => n1005, outb => n4018);
   U5042 : inv port map( inb => n1009, outb => n4021);
   U5043 : inv port map( inb => mult_125_G3_ab_3_7_port, outb => n1019);
   U5044 : inv port map( inb => n1037, outb => n4039);
   U5045 : inv port map( inb => n1041, outb => n4041);
   U5046 : inv port map( inb => mult_125_G3_ab_3_6_port, outb => n4044);
   U5047 : inv port map( inb => n1071, outb => n4058);
   U5048 : inv port map( inb => mult_125_G3_ab_3_5_port, outb => n1081);
   U5049 : inv port map( inb => n1104, outb => n4077);
   U5050 : inv port map( inb => mult_125_G3_ab_3_4_port, outb => n4080);
   U5051 : inv port map( inb => mult_125_G3_ab_3_3_port, outb => n1146);
   U5052 : inv port map( inb => mult_125_G3_ab_3_2_port, outb => n4115);
   U5053 : inv port map( inb => mult_125_G3_ab_3_1_port, outb => n4134);
   U5054 : inv port map( inb => n1208, outb => n4136);
   U5055 : inv port map( inb => n1237, outb => n4160);
   U5056 : inv port map( inb => n1241, outb => n4164);
   U5057 : inv port map( inb => n1245, outb => n4168);
   U5058 : inv port map( inb => n1249, outb => n4172);
   U5059 : inv port map( inb => n1253, outb => n4176);
   U5060 : inv port map( inb => mult_125_G2_ab_1_15_port, outb => n5211);
   U5061 : inv port map( inb => mult_125_G2_ab_2_14_port, outb => n5212);
   U5062 : inv port map( inb => n1284, outb => n4196);
   U5063 : inv port map( inb => n1288, outb => n4199);
   U5064 : inv port map( inb => n1292, outb => n4202);
   U5065 : inv port map( inb => n1296, outb => n4205);
   U5066 : inv port map( inb => n1300, outb => n4208);
   U5067 : inv port map( inb => mult_125_G2_ab_3_12_port, outb => n4211);
   U5068 : inv port map( inb => n1315, outb => n4218);
   U5069 : inv port map( inb => n1319, outb => n4221);
   U5070 : inv port map( inb => n1323, outb => n4224);
   U5071 : inv port map( inb => n1327, outb => n4227);
   U5072 : inv port map( inb => mult_125_G2_ab_3_11_port, outb => n1337);
   U5073 : inv port map( inb => n1347, outb => n4239);
   U5074 : inv port map( inb => n1351, outb => n4242);
   U5075 : inv port map( inb => n1355, outb => n4245);
   U5076 : inv port map( inb => n1359, outb => n4247);
   U5077 : inv port map( inb => mult_125_G2_ab_3_10_port, outb => n4250);
   U5078 : inv port map( inb => n1380, outb => n4259);
   U5079 : inv port map( inb => n1384, outb => n4262);
   U5080 : inv port map( inb => n1388, outb => n4265);
   U5081 : inv port map( inb => mult_125_G2_ab_3_9_port, outb => n4269);
   U5082 : inv port map( inb => n1411, outb => n4281);
   U5083 : inv port map( inb => n1415, outb => n4284);
   U5084 : inv port map( inb => n1419, outb => n4286);
   U5085 : inv port map( inb => mult_125_G2_ab_3_8_port, outb => n4289);
   U5086 : inv port map( inb => n1443, outb => n4303);
   U5087 : inv port map( inb => n1447, outb => n4306);
   U5088 : inv port map( inb => mult_125_G2_ab_3_7_port, outb => n1457);
   U5089 : inv port map( inb => n1475, outb => n4324);
   U5090 : inv port map( inb => n1479, outb => n4326);
   U5091 : inv port map( inb => mult_125_G2_ab_3_6_port, outb => n4329);
   U5092 : inv port map( inb => n1509, outb => n4343);
   U5093 : inv port map( inb => mult_125_G2_ab_3_5_port, outb => n1519);
   U5094 : inv port map( inb => n1542, outb => n4362);
   U5095 : inv port map( inb => mult_125_G2_ab_3_4_port, outb => n4365);
   U5096 : inv port map( inb => mult_125_G2_ab_3_3_port, outb => n1584);
   U5097 : inv port map( inb => mult_125_G2_ab_3_2_port, outb => n4400);
   U5098 : inv port map( inb => mult_125_G2_ab_3_1_port, outb => n4419);
   U5099 : inv port map( inb => n1646, outb => n4421);
   U5100 : inv port map( inb => n1675, outb => n4445);
   U5101 : inv port map( inb => n1679, outb => n4449);
   U5102 : inv port map( inb => n1683, outb => n4453);
   U5103 : inv port map( inb => n1687, outb => n4457);
   U5104 : inv port map( inb => n1691, outb => n4461);
   U5105 : inv port map( inb => mult_125_ab_1_15_port, outb => n5374);
   U5106 : inv port map( inb => mult_125_ab_2_14_port, outb => n5375);
   U5107 : inv port map( inb => n1722, outb => n4481);
   U5108 : inv port map( inb => n1726, outb => n4484);
   U5109 : inv port map( inb => n1730, outb => n4487);
   U5110 : inv port map( inb => n1734, outb => n4490);
   U5111 : inv port map( inb => n1738, outb => n4493);
   U5112 : inv port map( inb => mult_125_ab_3_12_port, outb => n4496);
   U5113 : inv port map( inb => n1753, outb => n4503);
   U5114 : inv port map( inb => n1757, outb => n4506);
   U5115 : inv port map( inb => n1761, outb => n4509);
   U5116 : inv port map( inb => n1765, outb => n4512);
   U5117 : inv port map( inb => mult_125_ab_3_11_port, outb => n1775);
   U5118 : inv port map( inb => n1785, outb => n4524);
   U5119 : inv port map( inb => n1789, outb => n4527);
   U5120 : inv port map( inb => n1793, outb => n4530);
   U5121 : inv port map( inb => n1797, outb => n4532);
   U5122 : inv port map( inb => mult_125_ab_3_10_port, outb => n4535);
   U5123 : inv port map( inb => n1818, outb => n4544);
   U5124 : inv port map( inb => n1822, outb => n4547);
   U5125 : inv port map( inb => n1826, outb => n4550);
   U5126 : inv port map( inb => mult_125_ab_3_9_port, outb => n4554);
   U5127 : inv port map( inb => n1849, outb => n4566);
   U5128 : inv port map( inb => n1853, outb => n4569);
   U5129 : inv port map( inb => n1857, outb => n4571);
   U5130 : inv port map( inb => mult_125_ab_3_8_port, outb => n4574);
   U5131 : inv port map( inb => n1881, outb => n4588);
   U5132 : inv port map( inb => n1885, outb => n4591);
   U5133 : inv port map( inb => mult_125_ab_3_7_port, outb => n1895);
   U5134 : inv port map( inb => n1913, outb => n4609);
   U5135 : inv port map( inb => n1917, outb => n4611);
   U5136 : inv port map( inb => mult_125_ab_3_6_port, outb => n4614);
   U5137 : inv port map( inb => n1947, outb => n4628);
   U5138 : inv port map( inb => mult_125_ab_3_5_port, outb => n1957);
   U5139 : inv port map( inb => n1980, outb => n4647);
   U5140 : inv port map( inb => mult_125_ab_3_4_port, outb => n4650);
   U5141 : inv port map( inb => mult_125_ab_3_3_port, outb => n2022);
   U5142 : inv port map( inb => mult_125_ab_3_2_port, outb => n4685);
   U5143 : inv port map( inb => mult_125_ab_3_1_port, outb => n4704);
   U5144 : inv port map( inb => n2084, outb => n4706);
   U5145 : inv port map( inb => n2113, outb => n4730);
   U5146 : inv port map( inb => n2117, outb => n4734);
   U5147 : inv port map( inb => n2121, outb => n4738);
   U5148 : inv port map( inb => n2125, outb => n4742);
   U5149 : inv port map( inb => n2129, outb => n4746);
   U5150 : inv port map( inb => mult_125_G4_ab_5_13_port, outb => n3624);
   U5151 : inv port map( inb => n4921, outb => n4924);
   U5152 : inv port map( inb => mult_125_G4_ab_7_11_port, outb => n3667);
   U5153 : inv port map( inb => mult_125_G4_ab_5_10_port, outb => n496);
   U5154 : inv port map( inb => mult_125_G4_ab_7_10_port, outb => n3685);
   U5155 : inv port map( inb => mult_125_G4_ab_9_9_port, outb => n3709);
   U5156 : inv port map( inb => mult_125_G4_ab_7_8_port, outb => n3726);
   U5157 : inv port map( inb => mult_125_G4_ab_9_8_port, outb => n3729);
   U5158 : inv port map( inb => mult_125_G4_ab_11_7_port, outb => n3752);
   U5159 : inv port map( inb => mult_125_G4_ab_9_6_port, outb => n625);
   U5160 : inv port map( inb => mult_125_G4_ab_11_6_port, outb => n3769);
   U5161 : inv port map( inb => mult_125_G4_ab_13_5_port, outb => n3791);
   U5162 : inv port map( inb => mult_125_G4_ab_11_4_port, outb => n693);
   U5163 : inv port map( inb => mult_125_G4_ab_13_4_port, outb => n3807);
   U5164 : inv port map( inb => mult_125_G3_ab_5_13_port, outb => n3909);
   U5165 : inv port map( inb => n5067, outb => n5070);
   U5166 : inv port map( inb => mult_125_G3_ab_7_11_port, outb => n3952);
   U5167 : inv port map( inb => mult_125_G3_ab_5_10_port, outb => n934);
   U5168 : inv port map( inb => mult_125_G3_ab_7_10_port, outb => n3970);
   U5169 : inv port map( inb => mult_125_G3_ab_9_9_port, outb => n3994);
   U5170 : inv port map( inb => mult_125_G3_ab_7_8_port, outb => n4011);
   U5171 : inv port map( inb => mult_125_G3_ab_9_8_port, outb => n4014);
   U5172 : inv port map( inb => mult_125_G3_ab_11_7_port, outb => n4037);
   U5173 : inv port map( inb => mult_125_G3_ab_9_6_port, outb => n1063);
   U5174 : inv port map( inb => mult_125_G3_ab_11_6_port, outb => n4054);
   U5175 : inv port map( inb => mult_125_G3_ab_13_5_port, outb => n4076);
   U5176 : inv port map( inb => mult_125_G3_ab_11_4_port, outb => n1131);
   U5177 : inv port map( inb => mult_125_G3_ab_13_4_port, outb => n4092);
   U5178 : inv port map( inb => mult_125_G2_ab_5_13_port, outb => n4194);
   U5179 : inv port map( inb => n5230, outb => n5233);
   U5180 : inv port map( inb => mult_125_G2_ab_7_11_port, outb => n4237);
   U5181 : inv port map( inb => mult_125_G2_ab_5_10_port, outb => n1372);
   U5182 : inv port map( inb => mult_125_G2_ab_7_10_port, outb => n4255);
   U5183 : inv port map( inb => mult_125_G2_ab_9_9_port, outb => n4279);
   U5184 : inv port map( inb => mult_125_G2_ab_7_8_port, outb => n4296);
   U5185 : inv port map( inb => mult_125_G2_ab_9_8_port, outb => n4299);
   U5186 : inv port map( inb => mult_125_G2_ab_11_7_port, outb => n4322);
   U5187 : inv port map( inb => mult_125_G2_ab_9_6_port, outb => n1501);
   U5188 : inv port map( inb => mult_125_G2_ab_11_6_port, outb => n4339);
   U5189 : inv port map( inb => mult_125_G2_ab_13_5_port, outb => n4361);
   U5190 : inv port map( inb => mult_125_G2_ab_11_4_port, outb => n1569);
   U5191 : inv port map( inb => mult_125_G2_ab_13_4_port, outb => n4377);
   U5192 : inv port map( inb => mult_125_ab_5_13_port, outb => n4479);
   U5193 : inv port map( inb => n5393, outb => n5396);
   U5194 : inv port map( inb => mult_125_ab_7_11_port, outb => n4522);
   U5195 : inv port map( inb => mult_125_ab_5_10_port, outb => n1810);
   U5196 : inv port map( inb => mult_125_ab_7_10_port, outb => n4540);
   U5197 : inv port map( inb => mult_125_ab_9_9_port, outb => n4564);
   U5198 : inv port map( inb => mult_125_ab_7_8_port, outb => n4581);
   U5199 : inv port map( inb => mult_125_ab_9_8_port, outb => n4584);
   U5200 : inv port map( inb => mult_125_ab_11_7_port, outb => n4607);
   U5201 : inv port map( inb => mult_125_ab_9_6_port, outb => n1939);
   U5202 : inv port map( inb => mult_125_ab_11_6_port, outb => n4624);
   U5203 : inv port map( inb => mult_125_ab_13_5_port, outb => n4646);
   U5204 : inv port map( inb => mult_125_ab_11_4_port, outb => n2007);
   U5205 : inv port map( inb => mult_125_ab_13_4_port, outb => n4662);
   U5206 : inv port map( inb => n4919, outb => n4922);
   U5207 : inv port map( inb => n396, outb => n4923);
   U5208 : inv port map( inb => n498, outb => n3684);
   U5209 : inv port map( inb => n561, outb => n3728);
   U5210 : inv port map( inb => n627, outb => n3768);
   U5211 : inv port map( inb => n695, outb => n3806);
   U5212 : inv port map( inb => n5065, outb => n5068);
   U5213 : inv port map( inb => n834, outb => n5069);
   U5214 : inv port map( inb => n936, outb => n3969);
   U5215 : inv port map( inb => n999, outb => n4013);
   U5216 : inv port map( inb => n1065, outb => n4053);
   U5217 : inv port map( inb => n1133, outb => n4091);
   U5218 : inv port map( inb => n5228, outb => n5231);
   U5219 : inv port map( inb => n1272, outb => n5232);
   U5220 : inv port map( inb => n1374, outb => n4254);
   U5221 : inv port map( inb => n1437, outb => n4298);
   U5222 : inv port map( inb => n1503, outb => n4338);
   U5223 : inv port map( inb => n1571, outb => n4376);
   U5224 : inv port map( inb => n5391, outb => n5394);
   U5225 : inv port map( inb => n1710, outb => n5395);
   U5226 : inv port map( inb => n1812, outb => n4539);
   U5227 : inv port map( inb => n1875, outb => n4583);
   U5228 : inv port map( inb => n1941, outb => n4623);
   U5229 : inv port map( inb => n2009, outb => n4661);
   U5230 : inv port map( inb => n400, outb => n3620);
   U5231 : inv port map( inb => n433, outb => n3643);
   U5232 : inv port map( inb => n470, outb => n3666);
   U5233 : inv port map( inb => n534, outb => n3708);
   U5234 : inv port map( inb => n598, outb => n3751);
   U5235 : inv port map( inb => n665, outb => n3790);
   U5236 : inv port map( inb => n703, outb => n4939);
   U5237 : inv port map( inb => n838, outb => n3905);
   U5238 : inv port map( inb => n871, outb => n3928);
   U5239 : inv port map( inb => n908, outb => n3951);
   U5240 : inv port map( inb => n972, outb => n3993);
   U5241 : inv port map( inb => n1036, outb => n4036);
   U5242 : inv port map( inb => n1103, outb => n4075);
   U5243 : inv port map( inb => n1141, outb => n5085);
   U5244 : inv port map( inb => n1276, outb => n4190);
   U5245 : inv port map( inb => n1309, outb => n4213);
   U5246 : inv port map( inb => n1346, outb => n4236);
   U5247 : inv port map( inb => n1410, outb => n4278);
   U5248 : inv port map( inb => n1474, outb => n4321);
   U5249 : inv port map( inb => n1541, outb => n4360);
   U5250 : inv port map( inb => n1579, outb => n5248);
   U5251 : inv port map( inb => n1714, outb => n4475);
   U5252 : inv port map( inb => n1747, outb => n4498);
   U5253 : inv port map( inb => n1784, outb => n4521);
   U5254 : inv port map( inb => n1848, outb => n4563);
   U5255 : inv port map( inb => n1912, outb => n4606);
   U5256 : inv port map( inb => n1979, outb => n4645);
   U5257 : inv port map( inb => n2017, outb => n5411);
   U5258 : inv port map( inb => mult_125_G4_ab_3_13_port, outb => n402);
   U5259 : inv port map( inb => n464, outb => n3661);
   U5260 : inv port map( inb => mult_125_G4_ab_4_11_port, outb => n3662);
   U5261 : inv port map( inb => mult_125_G4_ab_6_11_port, outb => n3665);
   U5262 : inv port map( inb => mult_125_G4_ab_6_9_port, outb => n3704);
   U5263 : inv port map( inb => n529, outb => n3706);
   U5264 : inv port map( inb => mult_125_G4_ab_8_9_port, outb => n3707);
   U5265 : inv port map( inb => mult_125_G4_ab_6_7_port, outb => n3744);
   U5266 : inv port map( inb => mult_125_G4_ab_8_7_port, outb => n3747);
   U5267 : inv port map( inb => n593, outb => n3749);
   U5268 : inv port map( inb => mult_125_G4_ab_10_7_port, outb => n3750);
   U5269 : inv port map( inb => mult_125_G4_ab_8_5_port, outb => n3783);
   U5270 : inv port map( inb => mult_125_G4_ab_10_5_port, outb => n3786);
   U5271 : inv port map( inb => n660, outb => n3788);
   U5272 : inv port map( inb => mult_125_G4_ab_12_5_port, outb => n3789);
   U5273 : inv port map( inb => n699, outb => n3808);
   U5274 : inv port map( inb => mult_125_G4_ab_10_3_port, outb => n3821);
   U5275 : inv port map( inb => mult_125_G4_ab_12_3_port, outb => n3824);
   U5276 : inv port map( inb => n728, outb => n3826);
   U5277 : inv port map( inb => mult_125_G4_ab_6_1_port, outb => n3854);
   U5278 : inv port map( inb => mult_125_G4_ab_8_1_port, outb => n3857);
   U5279 : inv port map( inb => mult_125_G4_ab_10_1_port, outb => n3860);
   U5280 : inv port map( inb => mult_125_G4_ab_12_1_port, outb => n3863);
   U5281 : inv port map( inb => mult_125_G3_ab_3_13_port, outb => n840);
   U5282 : inv port map( inb => n902, outb => n3946);
   U5283 : inv port map( inb => mult_125_G3_ab_4_11_port, outb => n3947);
   U5284 : inv port map( inb => mult_125_G3_ab_6_11_port, outb => n3950);
   U5285 : inv port map( inb => mult_125_G3_ab_6_9_port, outb => n3989);
   U5286 : inv port map( inb => n967, outb => n3991);
   U5287 : inv port map( inb => mult_125_G3_ab_8_9_port, outb => n3992);
   U5288 : inv port map( inb => mult_125_G3_ab_6_7_port, outb => n4029);
   U5289 : inv port map( inb => mult_125_G3_ab_8_7_port, outb => n4032);
   U5290 : inv port map( inb => n1031, outb => n4034);
   U5291 : inv port map( inb => mult_125_G3_ab_10_7_port, outb => n4035);
   U5292 : inv port map( inb => mult_125_G3_ab_8_5_port, outb => n4068);
   U5293 : inv port map( inb => mult_125_G3_ab_10_5_port, outb => n4071);
   U5294 : inv port map( inb => n1098, outb => n4073);
   U5295 : inv port map( inb => mult_125_G3_ab_12_5_port, outb => n4074);
   U5296 : inv port map( inb => n1137, outb => n4093);
   U5297 : inv port map( inb => mult_125_G3_ab_10_3_port, outb => n4106);
   U5298 : inv port map( inb => mult_125_G3_ab_12_3_port, outb => n4109);
   U5299 : inv port map( inb => n1166, outb => n4111);
   U5300 : inv port map( inb => mult_125_G3_ab_6_1_port, outb => n4139);
   U5301 : inv port map( inb => mult_125_G3_ab_8_1_port, outb => n4142);
   U5302 : inv port map( inb => mult_125_G3_ab_10_1_port, outb => n4145);
   U5303 : inv port map( inb => mult_125_G3_ab_12_1_port, outb => n4148);
   U5304 : inv port map( inb => mult_125_G2_ab_3_13_port, outb => n1278);
   U5305 : inv port map( inb => n1340, outb => n4231);
   U5306 : inv port map( inb => mult_125_G2_ab_4_11_port, outb => n4232);
   U5307 : inv port map( inb => mult_125_G2_ab_6_11_port, outb => n4235);
   U5308 : inv port map( inb => mult_125_G2_ab_6_9_port, outb => n4274);
   U5309 : inv port map( inb => n1405, outb => n4276);
   U5310 : inv port map( inb => mult_125_G2_ab_8_9_port, outb => n4277);
   U5311 : inv port map( inb => mult_125_G2_ab_6_7_port, outb => n4314);
   U5312 : inv port map( inb => mult_125_G2_ab_8_7_port, outb => n4317);
   U5313 : inv port map( inb => n1469, outb => n4319);
   U5314 : inv port map( inb => mult_125_G2_ab_10_7_port, outb => n4320);
   U5315 : inv port map( inb => mult_125_G2_ab_8_5_port, outb => n4353);
   U5316 : inv port map( inb => mult_125_G2_ab_10_5_port, outb => n4356);
   U5317 : inv port map( inb => n1536, outb => n4358);
   U5318 : inv port map( inb => mult_125_G2_ab_12_5_port, outb => n4359);
   U5319 : inv port map( inb => n1575, outb => n4378);
   U5320 : inv port map( inb => mult_125_G2_ab_10_3_port, outb => n4391);
   U5321 : inv port map( inb => mult_125_G2_ab_12_3_port, outb => n4394);
   U5322 : inv port map( inb => n1604, outb => n4396);
   U5323 : inv port map( inb => mult_125_G2_ab_6_1_port, outb => n4424);
   U5324 : inv port map( inb => mult_125_G2_ab_8_1_port, outb => n4427);
   U5325 : inv port map( inb => mult_125_G2_ab_10_1_port, outb => n4430);
   U5326 : inv port map( inb => mult_125_G2_ab_12_1_port, outb => n4433);
   U5327 : inv port map( inb => mult_125_ab_3_13_port, outb => n1716);
   U5328 : inv port map( inb => n1778, outb => n4516);
   U5329 : inv port map( inb => mult_125_ab_4_11_port, outb => n4517);
   U5330 : inv port map( inb => mult_125_ab_6_11_port, outb => n4520);
   U5331 : inv port map( inb => mult_125_ab_6_9_port, outb => n4559);
   U5332 : inv port map( inb => n1843, outb => n4561);
   U5333 : inv port map( inb => mult_125_ab_8_9_port, outb => n4562);
   U5334 : inv port map( inb => mult_125_ab_6_7_port, outb => n4599);
   U5335 : inv port map( inb => mult_125_ab_8_7_port, outb => n4602);
   U5336 : inv port map( inb => n1907, outb => n4604);
   U5337 : inv port map( inb => mult_125_ab_10_7_port, outb => n4605);
   U5338 : inv port map( inb => mult_125_ab_8_5_port, outb => n4638);
   U5339 : inv port map( inb => mult_125_ab_10_5_port, outb => n4641);
   U5340 : inv port map( inb => n1974, outb => n4643);
   U5341 : inv port map( inb => mult_125_ab_12_5_port, outb => n4644);
   U5342 : inv port map( inb => n2013, outb => n4663);
   U5343 : inv port map( inb => mult_125_ab_10_3_port, outb => n4676);
   U5344 : inv port map( inb => mult_125_ab_12_3_port, outb => n4679);
   U5345 : inv port map( inb => n2042, outb => n4681);
   U5346 : inv port map( inb => mult_125_ab_6_1_port, outb => n4709);
   U5347 : inv port map( inb => mult_125_ab_8_1_port, outb => n4712);
   U5348 : inv port map( inb => mult_125_ab_10_1_port, outb => n4715);
   U5349 : inv port map( inb => mult_125_ab_12_1_port, outb => n4718);
   U5350 : inv port map( inb => n3642, outb => n436);
   U5351 : inv port map( inb => n465, outb => n3664);
   U5352 : inv port map( inb => mult_125_G4_ab_13_2_port, outb => n3844);
   U5353 : inv port map( inb => n3927, outb => n874);
   U5354 : inv port map( inb => n903, outb => n3949);
   U5355 : inv port map( inb => mult_125_G3_ab_13_2_port, outb => n4129);
   U5356 : inv port map( inb => n4212, outb => n1312);
   U5357 : inv port map( inb => n1341, outb => n4234);
   U5358 : inv port map( inb => mult_125_G2_ab_13_2_port, outb => n4414);
   U5359 : inv port map( inb => n4497, outb => n1750);
   U5360 : inv port map( inb => n1779, outb => n4519);
   U5361 : inv port map( inb => mult_125_ab_13_2_port, outb => n4699);
   U5362 : inv port map( inb => n404, outb => n3623);
   U5363 : inv port map( inb => n493, outb => n3681);
   U5364 : inv port map( inb => n589, outb => n3746);
   U5365 : inv port map( inb => n656, outb => n3785);
   U5366 : inv port map( inb => n760, outb => n3846);
   U5367 : inv port map( inb => mult_125_G4_ab_15_2_port, outb => n4941);
   U5368 : inv port map( inb => n842, outb => n3908);
   U5369 : inv port map( inb => n931, outb => n3966);
   U5370 : inv port map( inb => n1027, outb => n4031);
   U5371 : inv port map( inb => n1094, outb => n4070);
   U5372 : inv port map( inb => n1198, outb => n4131);
   U5373 : inv port map( inb => mult_125_G3_ab_15_2_port, outb => n5087);
   U5374 : inv port map( inb => n1280, outb => n4193);
   U5375 : inv port map( inb => n1369, outb => n4251);
   U5376 : inv port map( inb => n1465, outb => n4316);
   U5377 : inv port map( inb => n1532, outb => n4355);
   U5378 : inv port map( inb => n1636, outb => n4416);
   U5379 : inv port map( inb => mult_125_G2_ab_15_2_port, outb => n5250);
   U5380 : inv port map( inb => n1718, outb => n4478);
   U5381 : inv port map( inb => n1807, outb => n4536);
   U5382 : inv port map( inb => n1903, outb => n4601);
   U5383 : inv port map( inb => n1970, outb => n4640);
   U5384 : inv port map( inb => n2074, outb => n4701);
   U5385 : inv port map( inb => mult_125_ab_15_2_port, outb => n5413);
   U5386 : inv port map( inb => mult_125_G4_ab_5_8_port, outb => n3723);
   U5387 : inv port map( inb => n557, outb => n3725);
   U5388 : inv port map( inb => mult_125_G4_ab_5_6_port, outb => n616);
   U5389 : inv port map( inb => mult_125_G4_ab_7_6_port, outb => n3764);
   U5390 : inv port map( inb => mult_125_G4_ab_5_4_port, outb => n679);
   U5391 : inv port map( inb => mult_125_G4_ab_7_4_port, outb => n684);
   U5392 : inv port map( inb => mult_125_G4_ab_9_4_port, outb => n3802);
   U5393 : inv port map( inb => mult_125_G4_ab_5_2_port, outb => n3833);
   U5394 : inv port map( inb => mult_125_G4_ab_7_2_port, outb => n746);
   U5395 : inv port map( inb => mult_125_G4_ab_9_2_port, outb => n3838);
   U5396 : inv port map( inb => mult_125_G4_ab_11_2_port, outb => n3841);
   U5397 : inv port map( inb => mult_125_G3_ab_5_8_port, outb => n4008);
   U5398 : inv port map( inb => n995, outb => n4010);
   U5399 : inv port map( inb => mult_125_G3_ab_5_6_port, outb => n1054);
   U5400 : inv port map( inb => mult_125_G3_ab_7_6_port, outb => n4049);
   U5401 : inv port map( inb => mult_125_G3_ab_5_4_port, outb => n1117);
   U5402 : inv port map( inb => mult_125_G3_ab_7_4_port, outb => n1122);
   U5403 : inv port map( inb => mult_125_G3_ab_9_4_port, outb => n4087);
   U5404 : inv port map( inb => mult_125_G3_ab_5_2_port, outb => n4118);
   U5405 : inv port map( inb => mult_125_G3_ab_7_2_port, outb => n1184);
   U5406 : inv port map( inb => mult_125_G3_ab_9_2_port, outb => n4123);
   U5407 : inv port map( inb => mult_125_G3_ab_11_2_port, outb => n4126);
   U5408 : inv port map( inb => mult_125_G2_ab_5_8_port, outb => n4293);
   U5409 : inv port map( inb => n1433, outb => n4295);
   U5410 : inv port map( inb => mult_125_G2_ab_5_6_port, outb => n1492);
   U5411 : inv port map( inb => mult_125_G2_ab_7_6_port, outb => n4334);
   U5412 : inv port map( inb => mult_125_G2_ab_5_4_port, outb => n1555);
   U5413 : inv port map( inb => mult_125_G2_ab_7_4_port, outb => n1560);
   U5414 : inv port map( inb => mult_125_G2_ab_9_4_port, outb => n4372);
   U5415 : inv port map( inb => mult_125_G2_ab_5_2_port, outb => n4403);
   U5416 : inv port map( inb => mult_125_G2_ab_7_2_port, outb => n1622);
   U5417 : inv port map( inb => mult_125_G2_ab_9_2_port, outb => n4408);
   U5418 : inv port map( inb => mult_125_G2_ab_11_2_port, outb => n4411);
   U5419 : inv port map( inb => mult_125_ab_5_8_port, outb => n4578);
   U5420 : inv port map( inb => n1871, outb => n4580);
   U5421 : inv port map( inb => mult_125_ab_5_6_port, outb => n1930);
   U5422 : inv port map( inb => mult_125_ab_7_6_port, outb => n4619);
   U5423 : inv port map( inb => mult_125_ab_5_4_port, outb => n1993);
   U5424 : inv port map( inb => mult_125_ab_7_4_port, outb => n1998);
   U5425 : inv port map( inb => mult_125_ab_9_4_port, outb => n4657);
   U5426 : inv port map( inb => mult_125_ab_5_2_port, outb => n4688);
   U5427 : inv port map( inb => mult_125_ab_7_2_port, outb => n2060);
   U5428 : inv port map( inb => mult_125_ab_9_2_port, outb => n4693);
   U5429 : inv port map( inb => mult_125_ab_11_2_port, outb => n4696);
   U5430 : inv port map( inb => n622, outb => n3765);
   U5431 : inv port map( inb => n686, outb => n3801);
   U5432 : inv port map( inb => n690, outb => n3803);
   U5433 : inv port map( inb => n732, outb => n4940);
   U5434 : inv port map( inb => n739, outb => n3832);
   U5435 : inv port map( inb => n748, outb => n3837);
   U5436 : inv port map( inb => n752, outb => n3840);
   U5437 : inv port map( inb => n756, outb => n3843);
   U5438 : inv port map( inb => n1060, outb => n4050);
   U5439 : inv port map( inb => n1124, outb => n4086);
   U5440 : inv port map( inb => n1128, outb => n4088);
   U5441 : inv port map( inb => n1170, outb => n5086);
   U5442 : inv port map( inb => n1177, outb => n4117);
   U5443 : inv port map( inb => n1186, outb => n4122);
   U5444 : inv port map( inb => n1190, outb => n4125);
   U5445 : inv port map( inb => n1194, outb => n4128);
   U5446 : inv port map( inb => n1498, outb => n4335);
   U5447 : inv port map( inb => n1562, outb => n4371);
   U5448 : inv port map( inb => n1566, outb => n4373);
   U5449 : inv port map( inb => n1608, outb => n5249);
   U5450 : inv port map( inb => n1615, outb => n4402);
   U5451 : inv port map( inb => n1624, outb => n4407);
   U5452 : inv port map( inb => n1628, outb => n4410);
   U5453 : inv port map( inb => n1632, outb => n4413);
   U5454 : inv port map( inb => n1936, outb => n4620);
   U5455 : inv port map( inb => n2000, outb => n4656);
   U5456 : inv port map( inb => n2004, outb => n4658);
   U5457 : inv port map( inb => n2046, outb => n5412);
   U5458 : inv port map( inb => n2053, outb => n4687);
   U5459 : inv port map( inb => n2062, outb => n4692);
   U5460 : inv port map( inb => n2066, outb => n4695);
   U5461 : inv port map( inb => n2070, outb => n4698);
   U5462 : inv port map( inb => n556, outb => n3722);
   U5463 : inv port map( inb => n618, outb => n3763);
   U5464 : inv port map( inb => n265, outb => mult_125_G4_A2_17_port);
   U5465 : inv port map( inb => n994, outb => n4007);
   U5466 : inv port map( inb => n1056, outb => n4048);
   U5467 : inv port map( inb => n373, outb => mult_125_G3_A2_17_port);
   U5468 : inv port map( inb => n1432, outb => n4292);
   U5469 : inv port map( inb => n1494, outb => n4333);
   U5470 : inv port map( inb => n337, outb => mult_125_G2_A2_17_port);
   U5471 : inv port map( inb => n1870, outb => n4577);
   U5472 : inv port map( inb => n1932, outb => n4618);
   U5473 : inv port map( inb => n301, outb => mult_125_A2_17_port);
   U5474 : inv port map( inb => n525, outb => n3703);
   U5475 : inv port map( inb => n584, outb => n3740);
   U5476 : inv port map( inb => mult_125_G4_ab_4_7_port, outb => n3741);
   U5477 : inv port map( inb => n585, outb => n3743);
   U5478 : inv port map( inb => mult_125_G4_ab_6_5_port, outb => n650);
   U5479 : inv port map( inb => n963, outb => n3988);
   U5480 : inv port map( inb => n1022, outb => n4025);
   U5481 : inv port map( inb => mult_125_G3_ab_4_7_port, outb => n4026);
   U5482 : inv port map( inb => n1023, outb => n4028);
   U5483 : inv port map( inb => mult_125_G3_ab_6_5_port, outb => n1088);
   U5484 : inv port map( inb => n1401, outb => n4273);
   U5485 : inv port map( inb => n1460, outb => n4310);
   U5486 : inv port map( inb => mult_125_G2_ab_4_7_port, outb => n4311);
   U5487 : inv port map( inb => n1461, outb => n4313);
   U5488 : inv port map( inb => mult_125_G2_ab_6_5_port, outb => n1526);
   U5489 : inv port map( inb => n1839, outb => n4558);
   U5490 : inv port map( inb => n1898, outb => n4595);
   U5491 : inv port map( inb => mult_125_ab_4_7_port, outb => n4596);
   U5492 : inv port map( inb => n1899, outb => n4598);
   U5493 : inv port map( inb => mult_125_ab_6_5_port, outb => n1964);
   U5494 : inv port map( inb => n524, outb => n3700);
   U5495 : inv port map( inb => mult_125_G4_ab_4_9_port, outb => n3701);
   U5496 : inv port map( inb => n652, outb => n3782);
   U5497 : inv port map( inb => n724, outb => n3823);
   U5498 : inv port map( inb => n962, outb => n3985);
   U5499 : inv port map( inb => mult_125_G3_ab_4_9_port, outb => n3986);
   U5500 : inv port map( inb => n1090, outb => n4067);
   U5501 : inv port map( inb => n1162, outb => n4108);
   U5502 : inv port map( inb => n1400, outb => n4270);
   U5503 : inv port map( inb => mult_125_G2_ab_4_9_port, outb => n4271);
   U5504 : inv port map( inb => n1528, outb => n4352);
   U5505 : inv port map( inb => n1600, outb => n4393);
   U5506 : inv port map( inb => n1838, outb => n4555);
   U5507 : inv port map( inb => mult_125_ab_4_9_port, outb => n4556);
   U5508 : inv port map( inb => n1966, outb => n4637);
   U5509 : inv port map( inb => n2038, outb => n4678);
   U5510 : inv port map( inb => mult_125_G4_ab_4_8_port, outb => n3721);
   U5511 : inv port map( inb => n681, outb => n3798);
   U5512 : inv port map( inb => n720, outb => n3820);
   U5513 : inv port map( inb => n743, outb => n3834);
   U5514 : inv port map( inb => mult_125_G3_ab_4_8_port, outb => n4006);
   U5515 : inv port map( inb => n1119, outb => n4083);
   U5516 : inv port map( inb => n1158, outb => n4105);
   U5517 : inv port map( inb => n1181, outb => n4119);
   U5518 : inv port map( inb => mult_125_G2_ab_4_8_port, outb => n4291);
   U5519 : inv port map( inb => n1557, outb => n4368);
   U5520 : inv port map( inb => n1596, outb => n4390);
   U5521 : inv port map( inb => n1619, outb => n4404);
   U5522 : inv port map( inb => mult_125_ab_4_8_port, outb => n4576);
   U5523 : inv port map( inb => n1995, outb => n4653);
   U5524 : inv port map( inb => n2034, outb => n4675);
   U5525 : inv port map( inb => n2057, outb => n4689);
   U5526 : inv port map( inb => n554, outb => n3720);
   U5527 : inv port map( inb => n646, outb => n3777);
   U5528 : inv port map( inb => mult_125_G4_ab_4_5_port, outb => n3778);
   U5529 : inv port map( inb => n711, outb => n3811);
   U5530 : inv port map( inb => mult_125_G4_ab_4_3_port, outb => n3812);
   U5531 : inv port map( inb => mult_125_G4_ab_6_3_port, outb => n3815);
   U5532 : inv port map( inb => mult_125_G4_ab_8_3_port, outb => n3818);
   U5533 : inv port map( inb => n992, outb => n4005);
   U5534 : inv port map( inb => n1084, outb => n4062);
   U5535 : inv port map( inb => mult_125_G3_ab_4_5_port, outb => n4063);
   U5536 : inv port map( inb => n1149, outb => n4096);
   U5537 : inv port map( inb => mult_125_G3_ab_4_3_port, outb => n4097);
   U5538 : inv port map( inb => mult_125_G3_ab_6_3_port, outb => n4100);
   U5539 : inv port map( inb => mult_125_G3_ab_8_3_port, outb => n4103);
   U5540 : inv port map( inb => n1430, outb => n4290);
   U5541 : inv port map( inb => n1522, outb => n4347);
   U5542 : inv port map( inb => mult_125_G2_ab_4_5_port, outb => n4348);
   U5543 : inv port map( inb => n1587, outb => n4381);
   U5544 : inv port map( inb => mult_125_G2_ab_4_3_port, outb => n4382);
   U5545 : inv port map( inb => mult_125_G2_ab_6_3_port, outb => n4385);
   U5546 : inv port map( inb => mult_125_G2_ab_8_3_port, outb => n4388);
   U5547 : inv port map( inb => n1868, outb => n4575);
   U5548 : inv port map( inb => n1960, outb => n4632);
   U5549 : inv port map( inb => mult_125_ab_4_5_port, outb => n4633);
   U5550 : inv port map( inb => n2025, outb => n4666);
   U5551 : inv port map( inb => mult_125_ab_4_3_port, outb => n4667);
   U5552 : inv port map( inb => mult_125_ab_6_3_port, outb => n4670);
   U5553 : inv port map( inb => mult_125_ab_8_3_port, outb => n4673);
   U5554 : inv port map( inb => n647, outb => n3779);
   U5555 : inv port map( inb => n716, outb => n3817);
   U5556 : inv port map( inb => n1085, outb => n4064);
   U5557 : inv port map( inb => n1154, outb => n4102);
   U5558 : inv port map( inb => n1523, outb => n4349);
   U5559 : inv port map( inb => n1592, outb => n4387);
   U5560 : inv port map( inb => n1961, outb => n4634);
   U5561 : inv port map( inb => n2030, outb => n4672);
   U5562 : inv port map( inb => n613, outb => n3760);
   U5563 : inv port map( inb => n676, outb => n3796);
   U5564 : inv port map( inb => n1051, outb => n4045);
   U5565 : inv port map( inb => n1114, outb => n4081);
   U5566 : inv port map( inb => n1489, outb => n4330);
   U5567 : inv port map( inb => n1552, outb => n4366);
   U5568 : inv port map( inb => n1927, outb => n4615);
   U5569 : inv port map( inb => n1990, outb => n4651);
   U5570 : inv port map( inb => n455, outb => n4927);
   U5571 : inv port map( inb => n516, outb => n4930);
   U5572 : inv port map( inb => n575, outb => n4933);
   U5573 : inv port map( inb => n637, outb => n4936);
   U5574 : inv port map( inb => n712, outb => n3814);
   U5575 : inv port map( inb => n775, outb => n3856);
   U5576 : inv port map( inb => n779, outb => n3859);
   U5577 : inv port map( inb => n783, outb => n3862);
   U5578 : inv port map( inb => n787, outb => n3865);
   U5579 : inv port map( inb => n791, outb => n4942);
   U5580 : inv port map( inb => n893, outb => n5073);
   U5581 : inv port map( inb => n954, outb => n5076);
   U5582 : inv port map( inb => n1013, outb => n5079);
   U5583 : inv port map( inb => n1075, outb => n5082);
   U5584 : inv port map( inb => n1150, outb => n4099);
   U5585 : inv port map( inb => n1213, outb => n4141);
   U5586 : inv port map( inb => n1217, outb => n4144);
   U5587 : inv port map( inb => n1221, outb => n4147);
   U5588 : inv port map( inb => n1225, outb => n4150);
   U5589 : inv port map( inb => n1229, outb => n5088);
   U5590 : inv port map( inb => n1331, outb => n5236);
   U5591 : inv port map( inb => n1392, outb => n5239);
   U5592 : inv port map( inb => n1451, outb => n5242);
   U5593 : inv port map( inb => n1513, outb => n5245);
   U5594 : inv port map( inb => n1588, outb => n4384);
   U5595 : inv port map( inb => n1651, outb => n4426);
   U5596 : inv port map( inb => n1655, outb => n4429);
   U5597 : inv port map( inb => n1659, outb => n4432);
   U5598 : inv port map( inb => n1663, outb => n4435);
   U5599 : inv port map( inb => n1667, outb => n5251);
   U5600 : inv port map( inb => n1769, outb => n5399);
   U5601 : inv port map( inb => n1830, outb => n5402);
   U5602 : inv port map( inb => n1889, outb => n5405);
   U5603 : inv port map( inb => n1951, outb => n5408);
   U5604 : inv port map( inb => n2026, outb => n4669);
   U5605 : inv port map( inb => n2089, outb => n4711);
   U5606 : inv port map( inb => n2093, outb => n4714);
   U5607 : inv port map( inb => n2097, outb => n4717);
   U5608 : inv port map( inb => n2101, outb => n4720);
   U5609 : inv port map( inb => n2105, outb => n5414);
   U5610 : inv port map( inb => n3625, outb => n411);
   U5611 : inv port map( inb => n3628, outb => n415);
   U5612 : inv port map( inb => n3631, outb => n419);
   U5613 : inv port map( inb => n3634, outb => n423);
   U5614 : inv port map( inb => mult_125_G4_ab_2_12_port, outb => n429);
   U5615 : inv port map( inb => n3639, outb => n432);
   U5616 : inv port map( inb => n3644, outb => n438);
   U5617 : inv port map( inb => n3647, outb => n442);
   U5618 : inv port map( inb => n3650, outb => n446);
   U5619 : inv port map( inb => n3653, outb => n450);
   U5620 : inv port map( inb => n3656, outb => n454);
   U5621 : inv port map( inb => mult_125_G4_ab_2_11_port, outb => n458);
   U5622 : inv port map( inb => n3668, outb => n474);
   U5623 : inv port map( inb => n3671, outb => n478);
   U5624 : inv port map( inb => n3674, outb => n482);
   U5625 : inv port map( inb => mult_125_G4_ab_15_11_port, outb => n486);
   U5626 : inv port map( inb => mult_125_G4_ab_2_10_port, outb => n489);
   U5627 : inv port map( inb => n3678, outb => n492);
   U5628 : inv port map( inb => n3688, outb => n507);
   U5629 : inv port map( inb => n3691, outb => n511);
   U5630 : inv port map( inb => n3694, outb => n515);
   U5631 : inv port map( inb => mult_125_G4_ab_2_9_port, outb => n519);
   U5632 : inv port map( inb => n3697, outb => n522);
   U5633 : inv port map( inb => n3705, outb => n532);
   U5634 : inv port map( inb => n3710, outb => n538);
   U5635 : inv port map( inb => n3713, outb => n542);
   U5636 : inv port map( inb => mult_125_G4_ab_15_9_port, outb => n546);
   U5637 : inv port map( inb => mult_125_G4_ab_2_8_port, outb => n549);
   U5638 : inv port map( inb => n3717, outb => n552);
   U5639 : inv port map( inb => n3724, outb => n560);
   U5640 : inv port map( inb => n3732, outb => n570);
   U5641 : inv port map( inb => n3735, outb => n574);
   U5642 : inv port map( inb => mult_125_G4_ab_2_7_port, outb => n578);
   U5643 : inv port map( inb => n3742, outb => n588);
   U5644 : inv port map( inb => n3745, outb => n592);
   U5645 : inv port map( inb => n3748, outb => n596);
   U5646 : inv port map( inb => n3753, outb => n602);
   U5647 : inv port map( inb => mult_125_G4_ab_15_7_port, outb => n606);
   U5648 : inv port map( inb => mult_125_G4_ab_2_6_port, outb => n609);
   U5649 : inv port map( inb => n3757, outb => n612);
   U5650 : inv port map( inb => n3762, outb => n621);
   U5651 : inv port map( inb => n3772, outb => n636);
   U5652 : inv port map( inb => mult_125_G4_ab_2_5_port, outb => n640);
   U5653 : inv port map( inb => n3784, outb => n659);
   U5654 : inv port map( inb => n3787, outb => n663);
   U5655 : inv port map( inb => mult_125_G4_ab_15_5_port, outb => n669);
   U5656 : inv port map( inb => mult_125_G4_ab_2_4_port, outb => n672);
   U5657 : inv port map( inb => n3793, outb => n675);
   U5658 : inv port map( inb => mult_125_G4_ab_15_4_port, outb => n702);
   U5659 : inv port map( inb => mult_125_G4_ab_2_3_port, outb => n705);
   U5660 : inv port map( inb => n3822, outb => n727);
   U5661 : inv port map( inb => mult_125_G4_ab_2_2_port, outb => n735);
   U5662 : inv port map( inb => n3828, outb => n738);
   U5663 : inv port map( inb => n3845, outb => n763);
   U5664 : inv port map( inb => mult_125_G4_ab_2_1_port, outb => n765);
   U5665 : inv port map( inb => n3847, outb => n768);
   U5666 : inv port map( inb => n771, outb => n3853);
   U5667 : inv port map( inb => n3855, outb => n778);
   U5668 : inv port map( inb => n3864, outb => n790);
   U5669 : inv port map( inb => n3874, outb => n802);
   U5670 : inv port map( inb => n3878, outb => n806);
   U5671 : inv port map( inb => n3882, outb => n810);
   U5672 : inv port map( inb => n3886, outb => n814);
   U5673 : inv port map( inb => n3890, outb => n818);
   U5674 : inv port map( inb => n821, outb => n240);
   U5675 : inv port map( inb => n3910, outb => n849);
   U5676 : inv port map( inb => n3913, outb => n853);
   U5677 : inv port map( inb => n3916, outb => n857);
   U5678 : inv port map( inb => n3919, outb => n861);
   U5679 : inv port map( inb => mult_125_G3_ab_2_12_port, outb => n867);
   U5680 : inv port map( inb => n3924, outb => n870);
   U5681 : inv port map( inb => n3929, outb => n876);
   U5682 : inv port map( inb => n3932, outb => n880);
   U5683 : inv port map( inb => n3935, outb => n884);
   U5684 : inv port map( inb => n3938, outb => n888);
   U5685 : inv port map( inb => n3941, outb => n892);
   U5686 : inv port map( inb => mult_125_G3_ab_2_11_port, outb => n896);
   U5687 : inv port map( inb => n3953, outb => n912);
   U5688 : inv port map( inb => n3956, outb => n916);
   U5689 : inv port map( inb => n3959, outb => n920);
   U5690 : inv port map( inb => mult_125_G3_ab_15_11_port, outb => n924);
   U5691 : inv port map( inb => mult_125_G3_ab_2_10_port, outb => n927);
   U5692 : inv port map( inb => n3963, outb => n930);
   U5693 : inv port map( inb => n3973, outb => n945);
   U5694 : inv port map( inb => n3976, outb => n949);
   U5695 : inv port map( inb => n3979, outb => n953);
   U5696 : inv port map( inb => mult_125_G3_ab_2_9_port, outb => n957);
   U5697 : inv port map( inb => n3982, outb => n960);
   U5698 : inv port map( inb => n3990, outb => n970);
   U5699 : inv port map( inb => n3995, outb => n976);
   U5700 : inv port map( inb => n3998, outb => n980);
   U5701 : inv port map( inb => mult_125_G3_ab_15_9_port, outb => n984);
   U5702 : inv port map( inb => mult_125_G3_ab_2_8_port, outb => n987);
   U5703 : inv port map( inb => n4002, outb => n990);
   U5704 : inv port map( inb => n4009, outb => n998);
   U5705 : inv port map( inb => n4017, outb => n1008);
   U5706 : inv port map( inb => n4020, outb => n1012);
   U5707 : inv port map( inb => mult_125_G3_ab_2_7_port, outb => n1016);
   U5708 : inv port map( inb => n4027, outb => n1026);
   U5709 : inv port map( inb => n4030, outb => n1030);
   U5710 : inv port map( inb => n4033, outb => n1034);
   U5711 : inv port map( inb => n4038, outb => n1040);
   U5712 : inv port map( inb => mult_125_G3_ab_15_7_port, outb => n1044);
   U5713 : inv port map( inb => mult_125_G3_ab_2_6_port, outb => n1047);
   U5714 : inv port map( inb => n4042, outb => n1050);
   U5715 : inv port map( inb => n4047, outb => n1059);
   U5716 : inv port map( inb => n4057, outb => n1074);
   U5717 : inv port map( inb => mult_125_G3_ab_2_5_port, outb => n1078);
   U5718 : inv port map( inb => n4069, outb => n1097);
   U5719 : inv port map( inb => n4072, outb => n1101);
   U5720 : inv port map( inb => mult_125_G3_ab_15_5_port, outb => n1107);
   U5721 : inv port map( inb => mult_125_G3_ab_2_4_port, outb => n1110);
   U5722 : inv port map( inb => n4078, outb => n1113);
   U5723 : inv port map( inb => mult_125_G3_ab_15_4_port, outb => n1140);
   U5724 : inv port map( inb => mult_125_G3_ab_2_3_port, outb => n1143);
   U5725 : inv port map( inb => n4107, outb => n1165);
   U5726 : inv port map( inb => mult_125_G3_ab_2_2_port, outb => n1173);
   U5727 : inv port map( inb => n4113, outb => n1176);
   U5728 : inv port map( inb => n4130, outb => n1201);
   U5729 : inv port map( inb => mult_125_G3_ab_2_1_port, outb => n1203);
   U5730 : inv port map( inb => n4132, outb => n1206);
   U5731 : inv port map( inb => n1209, outb => n4138);
   U5732 : inv port map( inb => n4140, outb => n1216);
   U5733 : inv port map( inb => n4149, outb => n1228);
   U5734 : inv port map( inb => n4159, outb => n1240);
   U5735 : inv port map( inb => n4163, outb => n1244);
   U5736 : inv port map( inb => n4167, outb => n1248);
   U5737 : inv port map( inb => n4171, outb => n1252);
   U5738 : inv port map( inb => n4175, outb => n1256);
   U5739 : inv port map( inb => n1259, outb => n348);
   U5740 : inv port map( inb => n4195, outb => n1287);
   U5741 : inv port map( inb => n4198, outb => n1291);
   U5742 : inv port map( inb => n4201, outb => n1295);
   U5743 : inv port map( inb => n4204, outb => n1299);
   U5744 : inv port map( inb => mult_125_G2_ab_2_12_port, outb => n1305);
   U5745 : inv port map( inb => n4209, outb => n1308);
   U5746 : inv port map( inb => n4214, outb => n1314);
   U5747 : inv port map( inb => n4217, outb => n1318);
   U5748 : inv port map( inb => n4220, outb => n1322);
   U5749 : inv port map( inb => n4223, outb => n1326);
   U5750 : inv port map( inb => n4226, outb => n1330);
   U5751 : inv port map( inb => mult_125_G2_ab_2_11_port, outb => n1334);
   U5752 : inv port map( inb => n4238, outb => n1350);
   U5753 : inv port map( inb => n4241, outb => n1354);
   U5754 : inv port map( inb => n4244, outb => n1358);
   U5755 : inv port map( inb => mult_125_G2_ab_15_11_port, outb => n1362);
   U5756 : inv port map( inb => mult_125_G2_ab_2_10_port, outb => n1365);
   U5757 : inv port map( inb => n4248, outb => n1368);
   U5758 : inv port map( inb => n4258, outb => n1383);
   U5759 : inv port map( inb => n4261, outb => n1387);
   U5760 : inv port map( inb => n4264, outb => n1391);
   U5761 : inv port map( inb => mult_125_G2_ab_2_9_port, outb => n1395);
   U5762 : inv port map( inb => n4267, outb => n1398);
   U5763 : inv port map( inb => n4275, outb => n1408);
   U5764 : inv port map( inb => n4280, outb => n1414);
   U5765 : inv port map( inb => n4283, outb => n1418);
   U5766 : inv port map( inb => mult_125_G2_ab_15_9_port, outb => n1422);
   U5767 : inv port map( inb => mult_125_G2_ab_2_8_port, outb => n1425);
   U5768 : inv port map( inb => n4287, outb => n1428);
   U5769 : inv port map( inb => n4294, outb => n1436);
   U5770 : inv port map( inb => n4302, outb => n1446);
   U5771 : inv port map( inb => n4305, outb => n1450);
   U5772 : inv port map( inb => mult_125_G2_ab_2_7_port, outb => n1454);
   U5773 : inv port map( inb => n4312, outb => n1464);
   U5774 : inv port map( inb => n4315, outb => n1468);
   U5775 : inv port map( inb => n4318, outb => n1472);
   U5776 : inv port map( inb => n4323, outb => n1478);
   U5777 : inv port map( inb => mult_125_G2_ab_15_7_port, outb => n1482);
   U5778 : inv port map( inb => mult_125_G2_ab_2_6_port, outb => n1485);
   U5779 : inv port map( inb => n4327, outb => n1488);
   U5780 : inv port map( inb => n4332, outb => n1497);
   U5781 : inv port map( inb => n4342, outb => n1512);
   U5782 : inv port map( inb => mult_125_G2_ab_2_5_port, outb => n1516);
   U5783 : inv port map( inb => n4354, outb => n1535);
   U5784 : inv port map( inb => n4357, outb => n1539);
   U5785 : inv port map( inb => mult_125_G2_ab_15_5_port, outb => n1545);
   U5786 : inv port map( inb => mult_125_G2_ab_2_4_port, outb => n1548);
   U5787 : inv port map( inb => n4363, outb => n1551);
   U5788 : inv port map( inb => mult_125_G2_ab_15_4_port, outb => n1578);
   U5789 : inv port map( inb => mult_125_G2_ab_2_3_port, outb => n1581);
   U5790 : inv port map( inb => n4392, outb => n1603);
   U5791 : inv port map( inb => mult_125_G2_ab_2_2_port, outb => n1611);
   U5792 : inv port map( inb => n4398, outb => n1614);
   U5793 : inv port map( inb => n4415, outb => n1639);
   U5794 : inv port map( inb => mult_125_G2_ab_2_1_port, outb => n1641);
   U5795 : inv port map( inb => n4417, outb => n1644);
   U5796 : inv port map( inb => n1647, outb => n4423);
   U5797 : inv port map( inb => n4425, outb => n1654);
   U5798 : inv port map( inb => n4434, outb => n1666);
   U5799 : inv port map( inb => n4444, outb => n1678);
   U5800 : inv port map( inb => n4448, outb => n1682);
   U5801 : inv port map( inb => n4452, outb => n1686);
   U5802 : inv port map( inb => n4456, outb => n1690);
   U5803 : inv port map( inb => n4460, outb => n1694);
   U5804 : inv port map( inb => n1697, outb => n312);
   U5805 : inv port map( inb => n4480, outb => n1725);
   U5806 : inv port map( inb => n4483, outb => n1729);
   U5807 : inv port map( inb => n4486, outb => n1733);
   U5808 : inv port map( inb => n4489, outb => n1737);
   U5809 : inv port map( inb => mult_125_ab_2_12_port, outb => n1743);
   U5810 : inv port map( inb => n4494, outb => n1746);
   U5811 : inv port map( inb => n4499, outb => n1752);
   U5812 : inv port map( inb => n4502, outb => n1756);
   U5813 : inv port map( inb => n4505, outb => n1760);
   U5814 : inv port map( inb => n4508, outb => n1764);
   U5815 : inv port map( inb => n4511, outb => n1768);
   U5816 : inv port map( inb => mult_125_ab_2_11_port, outb => n1772);
   U5817 : inv port map( inb => n4523, outb => n1788);
   U5818 : inv port map( inb => n4526, outb => n1792);
   U5819 : inv port map( inb => n4529, outb => n1796);
   U5820 : inv port map( inb => mult_125_ab_15_11_port, outb => n1800);
   U5821 : inv port map( inb => mult_125_ab_2_10_port, outb => n1803);
   U5822 : inv port map( inb => n4533, outb => n1806);
   U5823 : inv port map( inb => n4543, outb => n1821);
   U5824 : inv port map( inb => n4546, outb => n1825);
   U5825 : inv port map( inb => n4549, outb => n1829);
   U5826 : inv port map( inb => mult_125_ab_2_9_port, outb => n1833);
   U5827 : inv port map( inb => n4552, outb => n1836);
   U5828 : inv port map( inb => n4560, outb => n1846);
   U5829 : inv port map( inb => n4565, outb => n1852);
   U5830 : inv port map( inb => n4568, outb => n1856);
   U5831 : inv port map( inb => mult_125_ab_15_9_port, outb => n1860);
   U5832 : inv port map( inb => mult_125_ab_2_8_port, outb => n1863);
   U5833 : inv port map( inb => n4572, outb => n1866);
   U5834 : inv port map( inb => n4579, outb => n1874);
   U5835 : inv port map( inb => n4587, outb => n1884);
   U5836 : inv port map( inb => n4590, outb => n1888);
   U5837 : inv port map( inb => mult_125_ab_2_7_port, outb => n1892);
   U5838 : inv port map( inb => n4597, outb => n1902);
   U5839 : inv port map( inb => n4600, outb => n1906);
   U5840 : inv port map( inb => n4603, outb => n1910);
   U5841 : inv port map( inb => n4608, outb => n1916);
   U5842 : inv port map( inb => mult_125_ab_15_7_port, outb => n1920);
   U5843 : inv port map( inb => mult_125_ab_2_6_port, outb => n1923);
   U5844 : inv port map( inb => n4612, outb => n1926);
   U5845 : inv port map( inb => n4617, outb => n1935);
   U5846 : inv port map( inb => n4627, outb => n1950);
   U5847 : inv port map( inb => mult_125_ab_2_5_port, outb => n1954);
   U5848 : inv port map( inb => n4639, outb => n1973);
   U5849 : inv port map( inb => n4642, outb => n1977);
   U5850 : inv port map( inb => mult_125_ab_15_5_port, outb => n1983);
   U5851 : inv port map( inb => mult_125_ab_2_4_port, outb => n1986);
   U5852 : inv port map( inb => n4648, outb => n1989);
   U5853 : inv port map( inb => mult_125_ab_15_4_port, outb => n2016);
   U5854 : inv port map( inb => mult_125_ab_2_3_port, outb => n2019);
   U5855 : inv port map( inb => n4677, outb => n2041);
   U5856 : inv port map( inb => mult_125_ab_2_2_port, outb => n2049);
   U5857 : inv port map( inb => n4683, outb => n2052);
   U5858 : inv port map( inb => n4700, outb => n2077);
   U5859 : inv port map( inb => mult_125_ab_2_1_port, outb => n2079);
   U5860 : inv port map( inb => n4702, outb => n2082);
   U5861 : inv port map( inb => n2085, outb => n4708);
   U5862 : inv port map( inb => n4710, outb => n2092);
   U5863 : inv port map( inb => n4719, outb => n2104);
   U5864 : inv port map( inb => n4729, outb => n2116);
   U5865 : inv port map( inb => n4733, outb => n2120);
   U5866 : inv port map( inb => n4737, outb => n2124);
   U5867 : inv port map( inb => n4741, outb => n2128);
   U5868 : inv port map( inb => n4745, outb => n2132);
   U5869 : inv port map( inb => n2135, outb => n276);
   U5870 : inv port map( inb => multiplier_sigs_1_31_port, outb => n5270);
   U5871 : inv port map( inb => adder_mem_array_2_31_port, outb => n5269);
   U5872 : inv port map( inb => multiplier_sigs_0_31_port, outb => n5433);
   U5873 : inv port map( inb => adder_mem_array_1_31_port, outb => n5432);
   U5874 : inv port map( inb => multiplier_sigs_2_31_port, outb => n5107);
   U5875 : inv port map( inb => adder_mem_array_3_31_port, outb => n5106);
   U5876 : inv port map( inb => n2238, outb => n242);
   U5877 : inv port map( inb => mult_125_G4_ab_2_13_port, outb => n399);
   U5878 : inv port map( inb => n401, outb => n3621);
   U5879 : inv port map( inb => n3622, outb => n407);
   U5880 : inv port map( inb => n426, outb => n4926);
   U5881 : inv port map( inb => n435, outb => n3645);
   U5882 : inv port map( inb => n460, outb => n3660);
   U5883 : inv port map( inb => n3663, outb => n468);
   U5884 : inv port map( inb => n485, outb => n4929);
   U5885 : inv port map( inb => n4928, outb => n247);
   U5886 : inv port map( inb => mult_125_G4_ab_15_12_port, outb => n5037);
   U5887 : inv port map( inb => n495, outb => n3682);
   U5888 : inv port map( inb => n3683, outb => n501);
   U5889 : inv port map( inb => n3702, outb => n528);
   U5890 : inv port map( inb => n545, outb => n4932);
   U5891 : inv port map( inb => n4931, outb => n251);
   U5892 : inv port map( inb => mult_125_G4_ab_15_10_port, outb => n5038);
   U5893 : inv port map( inb => n3727, outb => n564);
   U5894 : inv port map( inb => n580, outb => n3739);
   U5895 : inv port map( inb => n605, outb => n4935);
   U5896 : inv port map( inb => n4934, outb => n255);
   U5897 : inv port map( inb => mult_125_G4_ab_15_8_port, outb => n5039);
   U5898 : inv port map( inb => n615, outb => n3761);
   U5899 : inv port map( inb => n624, outb => n3766);
   U5900 : inv port map( inb => n3767, outb => n630);
   U5901 : inv port map( inb => n642, outb => n3776);
   U5902 : inv port map( inb => n649, outb => n3780);
   U5903 : inv port map( inb => n3781, outb => n655);
   U5904 : inv port map( inb => n668, outb => n4938);
   U5905 : inv port map( inb => n4937, outb => n259);
   U5906 : inv port map( inb => mult_125_G4_ab_15_6_port, outb => n5040);
   U5907 : inv port map( inb => n678, outb => n3797);
   U5908 : inv port map( inb => n683, outb => n3799);
   U5909 : inv port map( inb => n3800, outb => n689);
   U5910 : inv port map( inb => n692, outb => n3804);
   U5911 : inv port map( inb => n3805, outb => n698);
   U5912 : inv port map( inb => n707, outb => n3810);
   U5913 : inv port map( inb => n3813, outb => n715);
   U5914 : inv port map( inb => n3816, outb => n719);
   U5915 : inv port map( inb => n3819, outb => n723);
   U5916 : inv port map( inb => n3825, outb => n731);
   U5917 : inv port map( inb => n3831, outb => n742);
   U5918 : inv port map( inb => n745, outb => n3835);
   U5919 : inv port map( inb => n3836, outb => n751);
   U5920 : inv port map( inb => n3839, outb => n755);
   U5921 : inv port map( inb => n3842, outb => n759);
   U5922 : inv port map( inb => n3852, outb => n774);
   U5923 : inv port map( inb => n3858, outb => n782);
   U5924 : inv port map( inb => n3861, outb => n786);
   U5925 : inv port map( inb => n793, outb => n3869);
   U5926 : inv port map( inb => n795, outb => n3871);
   U5927 : inv port map( inb => n3870, outb => n798);
   U5928 : inv port map( inb => n5041, outb => n5030);
   U5929 : inv port map( inb => mult_125_G4_ab_7_1_port, outb => n5042);
   U5930 : inv port map( inb => mult_125_G4_ab_9_1_port, outb => n5043);
   U5931 : inv port map( inb => mult_125_G4_ab_11_1_port, outb => n5044);
   U5932 : inv port map( inb => mult_125_G4_ab_13_1_port, outb => n5045);
   U5933 : inv port map( inb => mult_125_G4_ab_15_1_port, outb => n5046);
   U5934 : inv port map( inb => n2535, outb => n350);
   U5935 : inv port map( inb => mult_125_G3_ab_2_13_port, outb => n837);
   U5936 : inv port map( inb => n839, outb => n3906);
   U5937 : inv port map( inb => n3907, outb => n845);
   U5938 : inv port map( inb => n864, outb => n5072);
   U5939 : inv port map( inb => n873, outb => n3930);
   U5940 : inv port map( inb => n898, outb => n3945);
   U5941 : inv port map( inb => n3948, outb => n906);
   U5942 : inv port map( inb => n923, outb => n5075);
   U5943 : inv port map( inb => n5074, outb => n355);
   U5944 : inv port map( inb => mult_125_G3_ab_15_12_port, outb => n5200);
   U5945 : inv port map( inb => n933, outb => n3967);
   U5946 : inv port map( inb => n3968, outb => n939);
   U5947 : inv port map( inb => n3987, outb => n966);
   U5948 : inv port map( inb => n983, outb => n5078);
   U5949 : inv port map( inb => n5077, outb => n359);
   U5950 : inv port map( inb => mult_125_G3_ab_15_10_port, outb => n5201);
   U5951 : inv port map( inb => n4012, outb => n1002);
   U5952 : inv port map( inb => n1018, outb => n4024);
   U5953 : inv port map( inb => n1043, outb => n5081);
   U5954 : inv port map( inb => n5080, outb => n363);
   U5955 : inv port map( inb => mult_125_G3_ab_15_8_port, outb => n5202);
   U5956 : inv port map( inb => n1053, outb => n4046);
   U5957 : inv port map( inb => n1062, outb => n4051);
   U5958 : inv port map( inb => n4052, outb => n1068);
   U5959 : inv port map( inb => n1080, outb => n4061);
   U5960 : inv port map( inb => n1087, outb => n4065);
   U5961 : inv port map( inb => n4066, outb => n1093);
   U5962 : inv port map( inb => n1106, outb => n5084);
   U5963 : inv port map( inb => n5083, outb => n367);
   U5964 : inv port map( inb => mult_125_G3_ab_15_6_port, outb => n5203);
   U5965 : inv port map( inb => n1116, outb => n4082);
   U5966 : inv port map( inb => n1121, outb => n4084);
   U5967 : inv port map( inb => n4085, outb => n1127);
   U5968 : inv port map( inb => n1130, outb => n4089);
   U5969 : inv port map( inb => n4090, outb => n1136);
   U5970 : inv port map( inb => n1145, outb => n4095);
   U5971 : inv port map( inb => n4098, outb => n1153);
   U5972 : inv port map( inb => n4101, outb => n1157);
   U5973 : inv port map( inb => n4104, outb => n1161);
   U5974 : inv port map( inb => n4110, outb => n1169);
   U5975 : inv port map( inb => n4116, outb => n1180);
   U5976 : inv port map( inb => n1183, outb => n4120);
   U5977 : inv port map( inb => n4121, outb => n1189);
   U5978 : inv port map( inb => n4124, outb => n1193);
   U5979 : inv port map( inb => n4127, outb => n1197);
   U5980 : inv port map( inb => n4137, outb => n1212);
   U5981 : inv port map( inb => n4143, outb => n1220);
   U5982 : inv port map( inb => n4146, outb => n1224);
   U5983 : inv port map( inb => n1231, outb => n4154);
   U5984 : inv port map( inb => n1233, outb => n4156);
   U5985 : inv port map( inb => n4155, outb => n1236);
   U5986 : inv port map( inb => n5204, outb => n5193);
   U5987 : inv port map( inb => mult_125_G3_ab_7_1_port, outb => n5205);
   U5988 : inv port map( inb => mult_125_G3_ab_9_1_port, outb => n5206);
   U5989 : inv port map( inb => mult_125_G3_ab_11_1_port, outb => n5207);
   U5990 : inv port map( inb => mult_125_G3_ab_13_1_port, outb => n5208);
   U5991 : inv port map( inb => mult_125_G3_ab_15_1_port, outb => n5209);
   U5992 : inv port map( inb => n2832, outb => n314);
   U5993 : inv port map( inb => mult_125_G2_ab_2_13_port, outb => n1275);
   U5994 : inv port map( inb => n1277, outb => n4191);
   U5995 : inv port map( inb => n4192, outb => n1283);
   U5996 : inv port map( inb => n1302, outb => n5235);
   U5997 : inv port map( inb => n1311, outb => n4215);
   U5998 : inv port map( inb => n1336, outb => n4230);
   U5999 : inv port map( inb => n4233, outb => n1344);
   U6000 : inv port map( inb => n1361, outb => n5238);
   U6001 : inv port map( inb => n5237, outb => n319);
   U6002 : inv port map( inb => mult_125_G2_ab_15_12_port, outb => n5363);
   U6003 : inv port map( inb => n1371, outb => n4252);
   U6004 : inv port map( inb => n4253, outb => n1377);
   U6005 : inv port map( inb => n4272, outb => n1404);
   U6006 : inv port map( inb => n1421, outb => n5241);
   U6007 : inv port map( inb => n5240, outb => n323);
   U6008 : inv port map( inb => mult_125_G2_ab_15_10_port, outb => n5364);
   U6009 : inv port map( inb => n4297, outb => n1440);
   U6010 : inv port map( inb => n1456, outb => n4309);
   U6011 : inv port map( inb => n1481, outb => n5244);
   U6012 : inv port map( inb => n5243, outb => n327);
   U6013 : inv port map( inb => mult_125_G2_ab_15_8_port, outb => n5365);
   U6014 : inv port map( inb => n1491, outb => n4331);
   U6015 : inv port map( inb => n1500, outb => n4336);
   U6016 : inv port map( inb => n4337, outb => n1506);
   U6017 : inv port map( inb => n1518, outb => n4346);
   U6018 : inv port map( inb => n1525, outb => n4350);
   U6019 : inv port map( inb => n4351, outb => n1531);
   U6020 : inv port map( inb => n1544, outb => n5247);
   U6021 : inv port map( inb => n5246, outb => n331);
   U6022 : inv port map( inb => mult_125_G2_ab_15_6_port, outb => n5366);
   U6023 : inv port map( inb => n1554, outb => n4367);
   U6024 : inv port map( inb => n1559, outb => n4369);
   U6025 : inv port map( inb => n4370, outb => n1565);
   U6026 : inv port map( inb => n1568, outb => n4374);
   U6027 : inv port map( inb => n4375, outb => n1574);
   U6028 : inv port map( inb => n1583, outb => n4380);
   U6029 : inv port map( inb => n4383, outb => n1591);
   U6030 : inv port map( inb => n4386, outb => n1595);
   U6031 : inv port map( inb => n4389, outb => n1599);
   U6032 : inv port map( inb => n4395, outb => n1607);
   U6033 : inv port map( inb => n4401, outb => n1618);
   U6034 : inv port map( inb => n1621, outb => n4405);
   U6035 : inv port map( inb => n4406, outb => n1627);
   U6036 : inv port map( inb => n4409, outb => n1631);
   U6037 : inv port map( inb => n4412, outb => n1635);
   U6038 : inv port map( inb => n4422, outb => n1650);
   U6039 : inv port map( inb => n4428, outb => n1658);
   U6040 : inv port map( inb => n4431, outb => n1662);
   U6041 : inv port map( inb => n1669, outb => n4439);
   U6042 : inv port map( inb => n1671, outb => n4441);
   U6043 : inv port map( inb => n4440, outb => n1674);
   U6044 : inv port map( inb => n5367, outb => n5356);
   U6045 : inv port map( inb => mult_125_G2_ab_7_1_port, outb => n5368);
   U6046 : inv port map( inb => mult_125_G2_ab_9_1_port, outb => n5369);
   U6047 : inv port map( inb => mult_125_G2_ab_11_1_port, outb => n5370);
   U6048 : inv port map( inb => mult_125_G2_ab_13_1_port, outb => n5371);
   U6049 : inv port map( inb => mult_125_G2_ab_15_1_port, outb => n5372);
   U6050 : inv port map( inb => n3129, outb => n278);
   U6051 : inv port map( inb => mult_125_ab_2_13_port, outb => n1713);
   U6052 : inv port map( inb => n1715, outb => n4476);
   U6053 : inv port map( inb => n4477, outb => n1721);
   U6054 : inv port map( inb => n1740, outb => n5398);
   U6055 : inv port map( inb => n1749, outb => n4500);
   U6056 : inv port map( inb => n1774, outb => n4515);
   U6057 : inv port map( inb => n4518, outb => n1782);
   U6058 : inv port map( inb => n1799, outb => n5401);
   U6059 : inv port map( inb => n5400, outb => n283);
   U6060 : inv port map( inb => mult_125_ab_15_12_port, outb => n5526);
   U6061 : inv port map( inb => n1809, outb => n4537);
   U6062 : inv port map( inb => n4538, outb => n1815);
   U6063 : inv port map( inb => n4557, outb => n1842);
   U6064 : inv port map( inb => n1859, outb => n5404);
   U6065 : inv port map( inb => n5403, outb => n287);
   U6066 : inv port map( inb => mult_125_ab_15_10_port, outb => n5527);
   U6067 : inv port map( inb => n4582, outb => n1878);
   U6068 : inv port map( inb => n1894, outb => n4594);
   U6069 : inv port map( inb => n1919, outb => n5407);
   U6070 : inv port map( inb => n5406, outb => n291);
   U6071 : inv port map( inb => mult_125_ab_15_8_port, outb => n5528);
   U6072 : inv port map( inb => n1929, outb => n4616);
   U6073 : inv port map( inb => n1938, outb => n4621);
   U6074 : inv port map( inb => n4622, outb => n1944);
   U6075 : inv port map( inb => n1956, outb => n4631);
   U6076 : inv port map( inb => n1963, outb => n4635);
   U6077 : inv port map( inb => n4636, outb => n1969);
   U6078 : inv port map( inb => n1982, outb => n5410);
   U6079 : inv port map( inb => n5409, outb => n295);
   U6080 : inv port map( inb => mult_125_ab_15_6_port, outb => n5529);
   U6081 : inv port map( inb => n1992, outb => n4652);
   U6082 : inv port map( inb => n1997, outb => n4654);
   U6083 : inv port map( inb => n4655, outb => n2003);
   U6084 : inv port map( inb => n2006, outb => n4659);
   U6085 : inv port map( inb => n4660, outb => n2012);
   U6086 : inv port map( inb => n2021, outb => n4665);
   U6087 : inv port map( inb => n4668, outb => n2029);
   U6088 : inv port map( inb => n4671, outb => n2033);
   U6089 : inv port map( inb => n4674, outb => n2037);
   U6090 : inv port map( inb => n4680, outb => n2045);
   U6091 : inv port map( inb => n4686, outb => n2056);
   U6092 : inv port map( inb => n2059, outb => n4690);
   U6093 : inv port map( inb => n4691, outb => n2065);
   U6094 : inv port map( inb => n4694, outb => n2069);
   U6095 : inv port map( inb => n4697, outb => n2073);
   U6096 : inv port map( inb => n4707, outb => n2088);
   U6097 : inv port map( inb => n4713, outb => n2096);
   U6098 : inv port map( inb => n4716, outb => n2100);
   U6099 : inv port map( inb => n2107, outb => n4724);
   U6100 : inv port map( inb => n2109, outb => n4726);
   U6101 : inv port map( inb => n4725, outb => n2112);
   U6102 : inv port map( inb => n5530, outb => n5519);
   U6103 : inv port map( inb => mult_125_ab_7_1_port, outb => n5531);
   U6104 : inv port map( inb => mult_125_ab_9_1_port, outb => n5532);
   U6105 : inv port map( inb => mult_125_ab_11_1_port, outb => n5533);
   U6106 : inv port map( inb => mult_125_ab_13_1_port, outb => n5534);
   U6107 : inv port map( inb => mult_125_ab_15_1_port, outb => n5535);
   U6108 : inv port map( inb => n2136, outb => n5091);
   U6109 : inv port map( inb => n2163, outb => n5417);
   U6110 : inv port map( inb => n2166, outb => n5254);
   U6111 : inv port map( inb => n5536, outb => mult_125_G4_ZB);
   U6112 : inv port map( inb => n5537, outb => mult_125_G4_ZA);
   U6113 : inv port map( inb => n5538, outb => mult_125_G4_QB);
   U6114 : inv port map( inb => n5539, outb => mult_125_G4_QA);
   U6115 : inv port map( inb => mult_125_G4_A1_0_port, outb => n5540);
   U6116 : inv port map( inb => n5541, outb => multiplier_sigs_3_2_port);
   U6117 : inv port map( inb => mult_125_G4_A1_1_port, outb => n5542);
   U6118 : inv port map( inb => n5543, outb => multiplier_sigs_3_3_port);
   U6119 : inv port map( inb => mult_125_G4_A1_2_port, outb => n5544);
   U6120 : inv port map( inb => n5545, outb => multiplier_sigs_3_4_port);
   U6121 : inv port map( inb => mult_125_G4_A1_3_port, outb => n5546);
   U6122 : inv port map( inb => n5547, outb => multiplier_sigs_3_5_port);
   U6123 : inv port map( inb => mult_125_G4_A1_4_port, outb => n5548);
   U6124 : inv port map( inb => n5549, outb => multiplier_sigs_3_6_port);
   U6125 : inv port map( inb => mult_125_G4_A1_5_port, outb => n5550);
   U6126 : inv port map( inb => n5551, outb => multiplier_sigs_3_7_port);
   U6127 : inv port map( inb => mult_125_G4_A1_6_port, outb => n5552);
   U6128 : inv port map( inb => n5553, outb => multiplier_sigs_3_8_port);
   U6129 : inv port map( inb => mult_125_G4_A1_7_port, outb => n5554);
   U6130 : inv port map( inb => n5555, outb => multiplier_sigs_3_9_port);
   U6131 : inv port map( inb => mult_125_G4_A1_8_port, outb => n5556);
   U6132 : inv port map( inb => n5557, outb => multiplier_sigs_3_10_port);
   U6133 : inv port map( inb => mult_125_G4_A1_9_port, outb => n5558);
   U6134 : inv port map( inb => n5559, outb => multiplier_sigs_3_11_port);
   U6135 : inv port map( inb => mult_125_G4_A1_10_port, outb => n5560);
   U6136 : inv port map( inb => n5561, outb => multiplier_sigs_3_12_port);
   U6137 : inv port map( inb => mult_125_G4_A1_11_port, outb => n5562);
   U6138 : inv port map( inb => n5563, outb => multiplier_sigs_3_13_port);
   U6139 : inv port map( inb => mult_125_G4_A1_12_port, outb => n5564);
   U6140 : inv port map( inb => n5565, outb => multiplier_sigs_3_14_port);
   U6141 : inv port map( inb => mult_125_G4_A1_13_port, outb => n5566);
   U6142 : inv port map( inb => n5567, outb => multiplier_sigs_3_15_port);
   U6143 : inv port map( inb => mult_125_G4_A1_14_port, outb => n5568);
   U6144 : inv port map( inb => mult_125_G4_A2_14_port, outb => n5569);
   U6145 : inv port map( inb => n5570, outb => multiplier_sigs_3_16_port);
   U6146 : inv port map( inb => mult_125_G4_A1_15_port, outb => n5571);
   U6147 : inv port map( inb => mult_125_G4_A2_15_port, outb => n5572);
   U6148 : inv port map( inb => n5573, outb => 
                           mult_125_G4_FS_1_PG_int_0_3_3_port);
   U6149 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_3_2_port, outb => 
                           n5574);
   U6150 : inv port map( inb => mult_125_G4_FS_1_P_0_3_3_port, outb => n5575);
   U6151 : inv port map( inb => mult_125_G4_A1_16_port, outb => n5576);
   U6152 : inv port map( inb => mult_125_G4_A2_16_port, outb => n5577);
   U6153 : inv port map( inb => n5578, outb => 
                           mult_125_G4_FS_1_PG_int_0_4_0_port);
   U6154 : inv port map( inb => mult_125_G4_A1_17_port, outb => n5579);
   U6155 : inv port map( inb => mult_125_G4_A2_17_port, outb => n5580);
   U6156 : inv port map( inb => n5581, outb => 
                           mult_125_G4_FS_1_PG_int_0_4_1_port);
   U6157 : inv port map( inb => n5582, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_4_1_port);
   U6158 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_4_0_port, outb => 
                           n5583);
   U6159 : inv port map( inb => mult_125_G4_A1_18_port, outb => n5584);
   U6160 : inv port map( inb => mult_125_G4_A2_18_port, outb => n5585);
   U6161 : inv port map( inb => n5586, outb => 
                           mult_125_G4_FS_1_PG_int_0_4_2_port);
   U6162 : inv port map( inb => n5587, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_4_2_port);
   U6163 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_4_1_port, outb => 
                           n5588);
   U6164 : inv port map( inb => mult_125_G4_FS_1_C_1_4_1_port, outb => n5589);
   U6165 : inv port map( inb => mult_125_G4_FS_1_P_0_4_1_port, outb => n5590);
   U6166 : inv port map( inb => mult_125_G4_A1_19_port, outb => n5591);
   U6167 : inv port map( inb => mult_125_G4_A2_19_port, outb => n5592);
   U6168 : inv port map( inb => n5593, outb => 
                           mult_125_G4_FS_1_PG_int_0_4_3_port);
   U6169 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_4_2_port, outb => 
                           n5594);
   U6170 : inv port map( inb => mult_125_G4_FS_1_P_0_4_3_port, outb => n5595);
   U6171 : inv port map( inb => mult_125_G4_FS_1_C_1_4_2_port, outb => n5596);
   U6172 : inv port map( inb => mult_125_G4_FS_1_P_0_4_2_port, outb => n5597);
   U6173 : inv port map( inb => mult_125_G4_A1_20_port, outb => n5598);
   U6174 : inv port map( inb => mult_125_G4_A2_20_port, outb => n5599);
   U6175 : inv port map( inb => n5600, outb => 
                           mult_125_G4_FS_1_PG_int_0_5_0_port);
   U6176 : inv port map( inb => mult_125_G4_A1_21_port, outb => n5601);
   U6177 : inv port map( inb => mult_125_G4_A2_21_port, outb => n5602);
   U6178 : inv port map( inb => n5603, outb => 
                           mult_125_G4_FS_1_PG_int_0_5_1_port);
   U6179 : inv port map( inb => n5604, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_5_1_port);
   U6180 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_5_0_port, outb => 
                           n5605);
   U6181 : inv port map( inb => mult_125_G4_A1_22_port, outb => n5606);
   U6182 : inv port map( inb => mult_125_G4_A2_22_port, outb => n5607);
   U6183 : inv port map( inb => n5608, outb => 
                           mult_125_G4_FS_1_PG_int_0_5_2_port);
   U6184 : inv port map( inb => n5609, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_5_2_port);
   U6185 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_5_1_port, outb => 
                           n5610);
   U6186 : inv port map( inb => mult_125_G4_FS_1_C_1_5_1_port, outb => n5611);
   U6187 : inv port map( inb => mult_125_G4_FS_1_P_0_5_1_port, outb => n5612);
   U6188 : inv port map( inb => mult_125_G4_A1_23_port, outb => n5613);
   U6189 : inv port map( inb => mult_125_G4_A2_23_port, outb => n5614);
   U6190 : inv port map( inb => n5615, outb => 
                           mult_125_G4_FS_1_PG_int_0_5_3_port);
   U6191 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_5_2_port, outb => 
                           n5616);
   U6192 : inv port map( inb => mult_125_G4_FS_1_P_0_5_3_port, outb => n5617);
   U6193 : inv port map( inb => mult_125_G4_FS_1_C_1_5_2_port, outb => n5618);
   U6194 : inv port map( inb => mult_125_G4_FS_1_P_0_5_2_port, outb => n5619);
   U6195 : inv port map( inb => mult_125_G4_A1_24_port, outb => n5620);
   U6196 : inv port map( inb => mult_125_G4_A2_24_port, outb => n5621);
   U6197 : inv port map( inb => n5622, outb => 
                           mult_125_G4_FS_1_PG_int_0_6_0_port);
   U6198 : inv port map( inb => mult_125_G4_A1_25_port, outb => n5623);
   U6199 : inv port map( inb => mult_125_G4_A2_25_port, outb => n5624);
   U6200 : inv port map( inb => n5625, outb => 
                           mult_125_G4_FS_1_PG_int_0_6_1_port);
   U6201 : inv port map( inb => n5626, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_6_1_port);
   U6202 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_6_0_port, outb => 
                           n5627);
   U6203 : inv port map( inb => mult_125_G4_A1_26_port, outb => n5628);
   U6204 : inv port map( inb => mult_125_G4_A2_26_port, outb => n5629);
   U6205 : inv port map( inb => n5630, outb => 
                           mult_125_G4_FS_1_PG_int_0_6_2_port);
   U6206 : inv port map( inb => n5631, outb => 
                           mult_125_G4_FS_1_TEMP_P_0_6_2_port);
   U6207 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_6_1_port, outb => 
                           n5632);
   U6208 : inv port map( inb => mult_125_G4_FS_1_C_1_6_1_port, outb => n5633);
   U6209 : inv port map( inb => mult_125_G4_FS_1_P_0_6_1_port, outb => n5634);
   U6210 : inv port map( inb => mult_125_G4_A1_27_port, outb => n5635);
   U6211 : inv port map( inb => mult_125_G4_A2_27_port, outb => n5636);
   U6212 : inv port map( inb => n5637, outb => 
                           mult_125_G4_FS_1_PG_int_0_6_3_port);
   U6213 : inv port map( inb => mult_125_G4_FS_1_TEMP_G_0_6_2_port, outb => 
                           n5638);
   U6214 : inv port map( inb => mult_125_G4_FS_1_P_0_6_3_port, outb => n5639);
   U6215 : inv port map( inb => mult_125_G4_FS_1_C_1_6_2_port, outb => n5640);
   U6216 : inv port map( inb => mult_125_G4_FS_1_P_0_6_2_port, outb => n5641);
   U6217 : inv port map( inb => mult_125_G4_A1_28_port, outb => n5642);
   U6218 : inv port map( inb => mult_125_G4_A2_28_port, outb => n5643);
   U6219 : inv port map( inb => n5644, outb => 
                           mult_125_G4_FS_1_PG_int_0_7_0_port);
   U6220 : inv port map( inb => mult_125_G4_A1_29_port, outb => n5645);
   U6221 : inv port map( inb => mult_125_G4_A2_29_port, outb => n5646);
   U6222 : inv port map( inb => n5647, outb => 
                           mult_125_G4_FS_1_PG_int_0_7_1_port);
   U6223 : inv port map( inb => mult_125_G4_FS_1_C_1_7_0_port, outb => n5648);
   U6224 : inv port map( inb => mult_125_G4_FS_1_TEMP_P_0_7_0_port, outb => 
                           n5649);
   U6225 : inv port map( inb => mult_125_G4_FS_1_G_1_0_3_port, outb => n5650);
   U6226 : inv port map( inb => mult_125_G4_FS_1_C_1_4_0_port, outb => n5651);
   U6227 : inv port map( inb => mult_125_G4_FS_1_G_1_1_0_port, outb => n5653);
   U6228 : inv port map( inb => mult_125_G4_FS_1_C_1_5_0_port, outb => n5654);
   U6229 : inv port map( inb => mult_125_G4_FS_1_G_1_1_1_port, outb => n5656);
   U6230 : inv port map( inb => mult_125_G4_FS_1_C_1_6_0_port, outb => n5657);
   U6231 : inv port map( inb => mult_125_G4_FS_1_G_1_1_2_port, outb => n5659);
   U6232 : inv port map( inb => mult_125_G4_FS_1_G_2_0_0_port, outb => n5660);
   U6233 : inv port map( inb => n5661, outb => mult_125_ZB);
   U6234 : inv port map( inb => n5662, outb => mult_125_ZA);
   U6235 : inv port map( inb => n5663, outb => mult_125_QB);
   U6236 : inv port map( inb => n5664, outb => mult_125_QA);
   U6237 : inv port map( inb => mult_125_A1_0_port, outb => n5665);
   U6238 : inv port map( inb => n5666, outb => multiplier_sigs_0_2_port);
   U6239 : inv port map( inb => mult_125_A1_1_port, outb => n5667);
   U6240 : inv port map( inb => n5668, outb => multiplier_sigs_0_3_port);
   U6241 : inv port map( inb => mult_125_A1_2_port, outb => n5669);
   U6242 : inv port map( inb => n5670, outb => multiplier_sigs_0_4_port);
   U6243 : inv port map( inb => mult_125_A1_3_port, outb => n5671);
   U6244 : inv port map( inb => n5672, outb => multiplier_sigs_0_5_port);
   U6245 : inv port map( inb => mult_125_A1_4_port, outb => n5673);
   U6246 : inv port map( inb => n5674, outb => multiplier_sigs_0_6_port);
   U6247 : inv port map( inb => mult_125_A1_5_port, outb => n5675);
   U6248 : inv port map( inb => n5676, outb => multiplier_sigs_0_7_port);
   U6249 : inv port map( inb => mult_125_A1_6_port, outb => n5677);
   U6250 : inv port map( inb => n5678, outb => multiplier_sigs_0_8_port);
   U6251 : inv port map( inb => mult_125_A1_7_port, outb => n5679);
   U6252 : inv port map( inb => n5680, outb => multiplier_sigs_0_9_port);
   U6253 : inv port map( inb => mult_125_A1_8_port, outb => n5681);
   U6254 : inv port map( inb => n5682, outb => multiplier_sigs_0_10_port);
   U6255 : inv port map( inb => mult_125_A1_9_port, outb => n5683);
   U6256 : inv port map( inb => n5684, outb => multiplier_sigs_0_11_port);
   U6257 : inv port map( inb => mult_125_A1_10_port, outb => n5685);
   U6258 : inv port map( inb => n5686, outb => multiplier_sigs_0_12_port);
   U6259 : inv port map( inb => mult_125_A1_11_port, outb => n5687);
   U6260 : inv port map( inb => n5688, outb => multiplier_sigs_0_13_port);
   U6261 : inv port map( inb => mult_125_A1_12_port, outb => n5689);
   U6262 : inv port map( inb => n5690, outb => multiplier_sigs_0_14_port);
   U6263 : inv port map( inb => mult_125_A1_13_port, outb => n5691);
   U6264 : inv port map( inb => n5692, outb => multiplier_sigs_0_15_port);
   U6265 : inv port map( inb => mult_125_A1_14_port, outb => n5693);
   U6266 : inv port map( inb => mult_125_A2_14_port, outb => n5694);
   U6267 : inv port map( inb => n5695, outb => multiplier_sigs_0_16_port);
   U6268 : inv port map( inb => mult_125_A1_15_port, outb => n5696);
   U6269 : inv port map( inb => mult_125_A2_15_port, outb => n5697);
   U6270 : inv port map( inb => n5698, outb => mult_125_FS_1_PG_int_0_3_3_port)
                           ;
   U6271 : inv port map( inb => mult_125_FS_1_TEMP_G_0_3_2_port, outb => n5699)
                           ;
   U6272 : inv port map( inb => mult_125_FS_1_P_0_3_3_port, outb => n5700);
   U6273 : inv port map( inb => mult_125_A1_16_port, outb => n5701);
   U6274 : inv port map( inb => mult_125_A2_16_port, outb => n5702);
   U6275 : inv port map( inb => n5703, outb => mult_125_FS_1_PG_int_0_4_0_port)
                           ;
   U6276 : inv port map( inb => mult_125_A1_17_port, outb => n5704);
   U6277 : inv port map( inb => mult_125_A2_17_port, outb => n5705);
   U6278 : inv port map( inb => n5706, outb => mult_125_FS_1_PG_int_0_4_1_port)
                           ;
   U6279 : inv port map( inb => n5707, outb => mult_125_FS_1_TEMP_P_0_4_1_port)
                           ;
   U6280 : inv port map( inb => mult_125_FS_1_TEMP_P_0_4_0_port, outb => n5708)
                           ;
   U6281 : inv port map( inb => mult_125_A1_18_port, outb => n5709);
   U6282 : inv port map( inb => mult_125_A2_18_port, outb => n5710);
   U6283 : inv port map( inb => n5711, outb => mult_125_FS_1_PG_int_0_4_2_port)
                           ;
   U6284 : inv port map( inb => n5712, outb => mult_125_FS_1_TEMP_P_0_4_2_port)
                           ;
   U6285 : inv port map( inb => mult_125_FS_1_TEMP_G_0_4_1_port, outb => n5713)
                           ;
   U6286 : inv port map( inb => mult_125_FS_1_C_1_4_1_port, outb => n5714);
   U6287 : inv port map( inb => mult_125_FS_1_P_0_4_1_port, outb => n5715);
   U6288 : inv port map( inb => mult_125_A1_19_port, outb => n5716);
   U6289 : inv port map( inb => mult_125_A2_19_port, outb => n5717);
   U6290 : inv port map( inb => n5718, outb => mult_125_FS_1_PG_int_0_4_3_port)
                           ;
   U6291 : inv port map( inb => mult_125_FS_1_TEMP_G_0_4_2_port, outb => n5719)
                           ;
   U6292 : inv port map( inb => mult_125_FS_1_P_0_4_3_port, outb => n5720);
   U6293 : inv port map( inb => mult_125_FS_1_C_1_4_2_port, outb => n5721);
   U6294 : inv port map( inb => mult_125_FS_1_P_0_4_2_port, outb => n5722);
   U6295 : inv port map( inb => mult_125_A1_20_port, outb => n5723);
   U6296 : inv port map( inb => mult_125_A2_20_port, outb => n5724);
   U6297 : inv port map( inb => n5725, outb => mult_125_FS_1_PG_int_0_5_0_port)
                           ;
   U6298 : inv port map( inb => mult_125_A1_21_port, outb => n5726);
   U6299 : inv port map( inb => mult_125_A2_21_port, outb => n5727);
   U6300 : inv port map( inb => n5728, outb => mult_125_FS_1_PG_int_0_5_1_port)
                           ;
   U6301 : inv port map( inb => n5729, outb => mult_125_FS_1_TEMP_P_0_5_1_port)
                           ;
   U6302 : inv port map( inb => mult_125_FS_1_TEMP_P_0_5_0_port, outb => n5730)
                           ;
   U6303 : inv port map( inb => mult_125_A1_22_port, outb => n5731);
   U6304 : inv port map( inb => mult_125_A2_22_port, outb => n5732);
   U6305 : inv port map( inb => n5733, outb => mult_125_FS_1_PG_int_0_5_2_port)
                           ;
   U6306 : inv port map( inb => n5734, outb => mult_125_FS_1_TEMP_P_0_5_2_port)
                           ;
   U6307 : inv port map( inb => mult_125_FS_1_TEMP_G_0_5_1_port, outb => n5735)
                           ;
   U6308 : inv port map( inb => mult_125_FS_1_C_1_5_1_port, outb => n5736);
   U6309 : inv port map( inb => mult_125_FS_1_P_0_5_1_port, outb => n5737);
   U6310 : inv port map( inb => mult_125_A1_23_port, outb => n5738);
   U6311 : inv port map( inb => mult_125_A2_23_port, outb => n5739);
   U6312 : inv port map( inb => n5740, outb => mult_125_FS_1_PG_int_0_5_3_port)
                           ;
   U6313 : inv port map( inb => mult_125_FS_1_TEMP_G_0_5_2_port, outb => n5741)
                           ;
   U6314 : inv port map( inb => mult_125_FS_1_P_0_5_3_port, outb => n5742);
   U6315 : inv port map( inb => mult_125_FS_1_C_1_5_2_port, outb => n5743);
   U6316 : inv port map( inb => mult_125_FS_1_P_0_5_2_port, outb => n5744);
   U6317 : inv port map( inb => mult_125_A1_24_port, outb => n5745);
   U6318 : inv port map( inb => mult_125_A2_24_port, outb => n5746);
   U6319 : inv port map( inb => n5747, outb => mult_125_FS_1_PG_int_0_6_0_port)
                           ;
   U6320 : inv port map( inb => mult_125_A1_25_port, outb => n5748);
   U6321 : inv port map( inb => mult_125_A2_25_port, outb => n5749);
   U6322 : inv port map( inb => n5750, outb => mult_125_FS_1_PG_int_0_6_1_port)
                           ;
   U6323 : inv port map( inb => n5751, outb => mult_125_FS_1_TEMP_P_0_6_1_port)
                           ;
   U6324 : inv port map( inb => mult_125_FS_1_TEMP_P_0_6_0_port, outb => n5752)
                           ;
   U6325 : inv port map( inb => mult_125_A1_26_port, outb => n5753);
   U6326 : inv port map( inb => mult_125_A2_26_port, outb => n5754);
   U6327 : inv port map( inb => n5755, outb => mult_125_FS_1_PG_int_0_6_2_port)
                           ;
   U6328 : inv port map( inb => n5756, outb => mult_125_FS_1_TEMP_P_0_6_2_port)
                           ;
   U6329 : inv port map( inb => mult_125_FS_1_TEMP_G_0_6_1_port, outb => n5757)
                           ;
   U6330 : inv port map( inb => mult_125_FS_1_C_1_6_1_port, outb => n5758);
   U6331 : inv port map( inb => mult_125_FS_1_P_0_6_1_port, outb => n5759);
   U6332 : inv port map( inb => mult_125_A1_27_port, outb => n5760);
   U6333 : inv port map( inb => mult_125_A2_27_port, outb => n5761);
   U6334 : inv port map( inb => n5762, outb => mult_125_FS_1_PG_int_0_6_3_port)
                           ;
   U6335 : inv port map( inb => mult_125_FS_1_TEMP_G_0_6_2_port, outb => n5763)
                           ;
   U6336 : inv port map( inb => mult_125_FS_1_P_0_6_3_port, outb => n5764);
   U6337 : inv port map( inb => mult_125_FS_1_C_1_6_2_port, outb => n5765);
   U6338 : inv port map( inb => mult_125_FS_1_P_0_6_2_port, outb => n5766);
   U6339 : inv port map( inb => mult_125_A1_28_port, outb => n5767);
   U6340 : inv port map( inb => mult_125_A2_28_port, outb => n5768);
   U6341 : inv port map( inb => n5769, outb => mult_125_FS_1_PG_int_0_7_0_port)
                           ;
   U6342 : inv port map( inb => mult_125_A1_29_port, outb => n5770);
   U6343 : inv port map( inb => mult_125_A2_29_port, outb => n5771);
   U6344 : inv port map( inb => n5772, outb => mult_125_FS_1_PG_int_0_7_1_port)
                           ;
   U6345 : inv port map( inb => mult_125_FS_1_C_1_7_0_port, outb => n5773);
   U6346 : inv port map( inb => mult_125_FS_1_TEMP_P_0_7_0_port, outb => n5774)
                           ;
   U6347 : inv port map( inb => mult_125_FS_1_G_1_0_3_port, outb => n5775);
   U6348 : inv port map( inb => mult_125_FS_1_C_1_4_0_port, outb => n5776);
   U6349 : inv port map( inb => mult_125_FS_1_G_1_1_0_port, outb => n5778);
   U6350 : inv port map( inb => mult_125_FS_1_C_1_5_0_port, outb => n5779);
   U6351 : inv port map( inb => mult_125_FS_1_G_1_1_1_port, outb => n5781);
   U6352 : inv port map( inb => mult_125_FS_1_C_1_6_0_port, outb => n5782);
   U6353 : inv port map( inb => mult_125_FS_1_G_1_1_2_port, outb => n5784);
   U6354 : inv port map( inb => mult_125_FS_1_G_2_0_0_port, outb => n5785);
   U6355 : inv port map( inb => n5786, outb => mult_125_G2_ZB);
   U6356 : inv port map( inb => n5787, outb => mult_125_G2_ZA);
   U6357 : inv port map( inb => n5788, outb => mult_125_G2_QB);
   U6358 : inv port map( inb => n5789, outb => mult_125_G2_QA);
   U6359 : inv port map( inb => mult_125_G2_A1_0_port, outb => n5790);
   U6360 : inv port map( inb => n5791, outb => multiplier_sigs_1_2_port);
   U6361 : inv port map( inb => mult_125_G2_A1_1_port, outb => n5792);
   U6362 : inv port map( inb => n5793, outb => multiplier_sigs_1_3_port);
   U6363 : inv port map( inb => mult_125_G2_A1_2_port, outb => n5794);
   U6364 : inv port map( inb => n5795, outb => multiplier_sigs_1_4_port);
   U6365 : inv port map( inb => mult_125_G2_A1_3_port, outb => n5796);
   U6366 : inv port map( inb => n5797, outb => multiplier_sigs_1_5_port);
   U6367 : inv port map( inb => mult_125_G2_A1_4_port, outb => n5798);
   U6368 : inv port map( inb => n5799, outb => multiplier_sigs_1_6_port);
   U6369 : inv port map( inb => mult_125_G2_A1_5_port, outb => n5800);
   U6370 : inv port map( inb => n5801, outb => multiplier_sigs_1_7_port);
   U6371 : inv port map( inb => mult_125_G2_A1_6_port, outb => n5802);
   U6372 : inv port map( inb => n5803, outb => multiplier_sigs_1_8_port);
   U6373 : inv port map( inb => mult_125_G2_A1_7_port, outb => n5804);
   U6374 : inv port map( inb => n5805, outb => multiplier_sigs_1_9_port);
   U6375 : inv port map( inb => mult_125_G2_A1_8_port, outb => n5806);
   U6376 : inv port map( inb => n5807, outb => multiplier_sigs_1_10_port);
   U6377 : inv port map( inb => mult_125_G2_A1_9_port, outb => n5808);
   U6378 : inv port map( inb => n5809, outb => multiplier_sigs_1_11_port);
   U6379 : inv port map( inb => mult_125_G2_A1_10_port, outb => n5810);
   U6380 : inv port map( inb => n5811, outb => multiplier_sigs_1_12_port);
   U6381 : inv port map( inb => mult_125_G2_A1_11_port, outb => n5812);
   U6382 : inv port map( inb => n5813, outb => multiplier_sigs_1_13_port);
   U6383 : inv port map( inb => mult_125_G2_A1_12_port, outb => n5814);
   U6384 : inv port map( inb => n5815, outb => multiplier_sigs_1_14_port);
   U6385 : inv port map( inb => mult_125_G2_A1_13_port, outb => n5816);
   U6386 : inv port map( inb => n5817, outb => multiplier_sigs_1_15_port);
   U6387 : inv port map( inb => mult_125_G2_A1_14_port, outb => n5818);
   U6388 : inv port map( inb => mult_125_G2_A2_14_port, outb => n5819);
   U6389 : inv port map( inb => n5820, outb => multiplier_sigs_1_16_port);
   U6390 : inv port map( inb => mult_125_G2_A1_15_port, outb => n5821);
   U6391 : inv port map( inb => mult_125_G2_A2_15_port, outb => n5822);
   U6392 : inv port map( inb => n5823, outb => 
                           mult_125_G2_FS_1_PG_int_0_3_3_port);
   U6393 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_3_2_port, outb => 
                           n5824);
   U6394 : inv port map( inb => mult_125_G2_FS_1_P_0_3_3_port, outb => n5825);
   U6395 : inv port map( inb => mult_125_G2_A1_16_port, outb => n5826);
   U6396 : inv port map( inb => mult_125_G2_A2_16_port, outb => n5827);
   U6397 : inv port map( inb => n5828, outb => 
                           mult_125_G2_FS_1_PG_int_0_4_0_port);
   U6398 : inv port map( inb => mult_125_G2_A1_17_port, outb => n5829);
   U6399 : inv port map( inb => mult_125_G2_A2_17_port, outb => n5830);
   U6400 : inv port map( inb => n5831, outb => 
                           mult_125_G2_FS_1_PG_int_0_4_1_port);
   U6401 : inv port map( inb => n5832, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_4_1_port);
   U6402 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_4_0_port, outb => 
                           n5833);
   U6403 : inv port map( inb => mult_125_G2_A1_18_port, outb => n5834);
   U6404 : inv port map( inb => mult_125_G2_A2_18_port, outb => n5835);
   U6405 : inv port map( inb => n5836, outb => 
                           mult_125_G2_FS_1_PG_int_0_4_2_port);
   U6406 : inv port map( inb => n5837, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_4_2_port);
   U6407 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_4_1_port, outb => 
                           n5838);
   U6408 : inv port map( inb => mult_125_G2_FS_1_C_1_4_1_port, outb => n5839);
   U6409 : inv port map( inb => mult_125_G2_FS_1_P_0_4_1_port, outb => n5840);
   U6410 : inv port map( inb => mult_125_G2_A1_19_port, outb => n5841);
   U6411 : inv port map( inb => mult_125_G2_A2_19_port, outb => n5842);
   U6412 : inv port map( inb => n5843, outb => 
                           mult_125_G2_FS_1_PG_int_0_4_3_port);
   U6413 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_4_2_port, outb => 
                           n5844);
   U6414 : inv port map( inb => mult_125_G2_FS_1_P_0_4_3_port, outb => n5845);
   U6415 : inv port map( inb => mult_125_G2_FS_1_C_1_4_2_port, outb => n5846);
   U6416 : inv port map( inb => mult_125_G2_FS_1_P_0_4_2_port, outb => n5847);
   U6417 : inv port map( inb => mult_125_G2_A1_20_port, outb => n5848);
   U6418 : inv port map( inb => mult_125_G2_A2_20_port, outb => n5849);
   U6419 : inv port map( inb => n5850, outb => 
                           mult_125_G2_FS_1_PG_int_0_5_0_port);
   U6420 : inv port map( inb => mult_125_G2_A1_21_port, outb => n5851);
   U6421 : inv port map( inb => mult_125_G2_A2_21_port, outb => n5852);
   U6422 : inv port map( inb => n5853, outb => 
                           mult_125_G2_FS_1_PG_int_0_5_1_port);
   U6423 : inv port map( inb => n5854, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_5_1_port);
   U6424 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_5_0_port, outb => 
                           n5855);
   U6425 : inv port map( inb => mult_125_G2_A1_22_port, outb => n5856);
   U6426 : inv port map( inb => mult_125_G2_A2_22_port, outb => n5857);
   U6427 : inv port map( inb => n5858, outb => 
                           mult_125_G2_FS_1_PG_int_0_5_2_port);
   U6428 : inv port map( inb => n5859, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_5_2_port);
   U6429 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_5_1_port, outb => 
                           n5860);
   U6430 : inv port map( inb => mult_125_G2_FS_1_C_1_5_1_port, outb => n5861);
   U6431 : inv port map( inb => mult_125_G2_FS_1_P_0_5_1_port, outb => n5862);
   U6432 : inv port map( inb => mult_125_G2_A1_23_port, outb => n5863);
   U6433 : inv port map( inb => mult_125_G2_A2_23_port, outb => n5864);
   U6434 : inv port map( inb => n5865, outb => 
                           mult_125_G2_FS_1_PG_int_0_5_3_port);
   U6435 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_5_2_port, outb => 
                           n5866);
   U6436 : inv port map( inb => mult_125_G2_FS_1_P_0_5_3_port, outb => n5867);
   U6437 : inv port map( inb => mult_125_G2_FS_1_C_1_5_2_port, outb => n5868);
   U6438 : inv port map( inb => mult_125_G2_FS_1_P_0_5_2_port, outb => n5869);
   U6439 : inv port map( inb => mult_125_G2_A1_24_port, outb => n5870);
   U6440 : inv port map( inb => mult_125_G2_A2_24_port, outb => n5871);
   U6441 : inv port map( inb => n5872, outb => 
                           mult_125_G2_FS_1_PG_int_0_6_0_port);
   U6442 : inv port map( inb => mult_125_G2_A1_25_port, outb => n5873);
   U6443 : inv port map( inb => mult_125_G2_A2_25_port, outb => n5874);
   U6444 : inv port map( inb => n5875, outb => 
                           mult_125_G2_FS_1_PG_int_0_6_1_port);
   U6445 : inv port map( inb => n5876, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_6_1_port);
   U6446 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_6_0_port, outb => 
                           n5877);
   U6447 : inv port map( inb => mult_125_G2_A1_26_port, outb => n5878);
   U6448 : inv port map( inb => mult_125_G2_A2_26_port, outb => n5879);
   U6449 : inv port map( inb => n5880, outb => 
                           mult_125_G2_FS_1_PG_int_0_6_2_port);
   U6450 : inv port map( inb => n5881, outb => 
                           mult_125_G2_FS_1_TEMP_P_0_6_2_port);
   U6451 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_6_1_port, outb => 
                           n5882);
   U6452 : inv port map( inb => mult_125_G2_FS_1_C_1_6_1_port, outb => n5883);
   U6453 : inv port map( inb => mult_125_G2_FS_1_P_0_6_1_port, outb => n5884);
   U6454 : inv port map( inb => mult_125_G2_A1_27_port, outb => n5885);
   U6455 : inv port map( inb => mult_125_G2_A2_27_port, outb => n5886);
   U6456 : inv port map( inb => n5887, outb => 
                           mult_125_G2_FS_1_PG_int_0_6_3_port);
   U6457 : inv port map( inb => mult_125_G2_FS_1_TEMP_G_0_6_2_port, outb => 
                           n5888);
   U6458 : inv port map( inb => mult_125_G2_FS_1_P_0_6_3_port, outb => n5889);
   U6459 : inv port map( inb => mult_125_G2_FS_1_C_1_6_2_port, outb => n5890);
   U6460 : inv port map( inb => mult_125_G2_FS_1_P_0_6_2_port, outb => n5891);
   U6461 : inv port map( inb => mult_125_G2_A1_28_port, outb => n5892);
   U6462 : inv port map( inb => mult_125_G2_A2_28_port, outb => n5893);
   U6463 : inv port map( inb => n5894, outb => 
                           mult_125_G2_FS_1_PG_int_0_7_0_port);
   U6464 : inv port map( inb => mult_125_G2_A1_29_port, outb => n5895);
   U6465 : inv port map( inb => mult_125_G2_A2_29_port, outb => n5896);
   U6466 : inv port map( inb => n5897, outb => 
                           mult_125_G2_FS_1_PG_int_0_7_1_port);
   U6467 : inv port map( inb => mult_125_G2_FS_1_C_1_7_0_port, outb => n5898);
   U6468 : inv port map( inb => mult_125_G2_FS_1_TEMP_P_0_7_0_port, outb => 
                           n5899);
   U6469 : inv port map( inb => mult_125_G2_FS_1_G_1_0_3_port, outb => n5900);
   U6470 : inv port map( inb => mult_125_G2_FS_1_C_1_4_0_port, outb => n5901);
   U6471 : inv port map( inb => mult_125_G2_FS_1_G_1_1_0_port, outb => n5903);
   U6472 : inv port map( inb => mult_125_G2_FS_1_C_1_5_0_port, outb => n5904);
   U6473 : inv port map( inb => mult_125_G2_FS_1_G_1_1_1_port, outb => n5906);
   U6474 : inv port map( inb => mult_125_G2_FS_1_C_1_6_0_port, outb => n5907);
   U6475 : inv port map( inb => mult_125_G2_FS_1_G_1_1_2_port, outb => n5909);
   U6476 : inv port map( inb => mult_125_G2_FS_1_G_2_0_0_port, outb => n5910);
   U6477 : inv port map( inb => n5911, outb => mult_125_G3_ZB);
   U6478 : inv port map( inb => n5912, outb => mult_125_G3_ZA);
   U6479 : inv port map( inb => n5913, outb => mult_125_G3_QB);
   U6480 : inv port map( inb => n5914, outb => mult_125_G3_QA);
   U6481 : inv port map( inb => mult_125_G3_A1_0_port, outb => n5915);
   U6482 : inv port map( inb => n5916, outb => multiplier_sigs_2_2_port);
   U6483 : inv port map( inb => mult_125_G3_A1_1_port, outb => n5917);
   U6484 : inv port map( inb => n5918, outb => multiplier_sigs_2_3_port);
   U6485 : inv port map( inb => mult_125_G3_A1_2_port, outb => n5919);
   U6486 : inv port map( inb => n5920, outb => multiplier_sigs_2_4_port);
   U6487 : inv port map( inb => mult_125_G3_A1_3_port, outb => n5921);
   U6488 : inv port map( inb => n5922, outb => multiplier_sigs_2_5_port);
   U6489 : inv port map( inb => mult_125_G3_A1_4_port, outb => n5923);
   U6490 : inv port map( inb => n5924, outb => multiplier_sigs_2_6_port);
   U6491 : inv port map( inb => mult_125_G3_A1_5_port, outb => n5925);
   U6492 : inv port map( inb => n5926, outb => multiplier_sigs_2_7_port);
   U6493 : inv port map( inb => mult_125_G3_A1_6_port, outb => n5927);
   U6494 : inv port map( inb => n5928, outb => multiplier_sigs_2_8_port);
   U6495 : inv port map( inb => mult_125_G3_A1_7_port, outb => n5929);
   U6496 : inv port map( inb => n5930, outb => multiplier_sigs_2_9_port);
   U6497 : inv port map( inb => mult_125_G3_A1_8_port, outb => n5931);
   U6498 : inv port map( inb => n5932, outb => multiplier_sigs_2_10_port);
   U6499 : inv port map( inb => mult_125_G3_A1_9_port, outb => n5933);
   U6500 : inv port map( inb => n5934, outb => multiplier_sigs_2_11_port);
   U6501 : inv port map( inb => mult_125_G3_A1_10_port, outb => n5935);
   U6502 : inv port map( inb => n5936, outb => multiplier_sigs_2_12_port);
   U6503 : inv port map( inb => mult_125_G3_A1_11_port, outb => n5937);
   U6504 : inv port map( inb => n5938, outb => multiplier_sigs_2_13_port);
   U6505 : inv port map( inb => mult_125_G3_A1_12_port, outb => n5939);
   U6506 : inv port map( inb => n5940, outb => multiplier_sigs_2_14_port);
   U6507 : inv port map( inb => mult_125_G3_A1_13_port, outb => n5941);
   U6508 : inv port map( inb => n5942, outb => multiplier_sigs_2_15_port);
   U6509 : inv port map( inb => mult_125_G3_A1_14_port, outb => n5943);
   U6510 : inv port map( inb => mult_125_G3_A2_14_port, outb => n5944);
   U6511 : inv port map( inb => n5945, outb => multiplier_sigs_2_16_port);
   U6512 : inv port map( inb => mult_125_G3_A1_15_port, outb => n5946);
   U6513 : inv port map( inb => mult_125_G3_A2_15_port, outb => n5947);
   U6514 : inv port map( inb => n5948, outb => 
                           mult_125_G3_FS_1_PG_int_0_3_3_port);
   U6515 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_3_2_port, outb => 
                           n5949);
   U6516 : inv port map( inb => mult_125_G3_FS_1_P_0_3_3_port, outb => n5950);
   U6517 : inv port map( inb => mult_125_G3_A1_16_port, outb => n5951);
   U6518 : inv port map( inb => mult_125_G3_A2_16_port, outb => n5952);
   U6519 : inv port map( inb => n5953, outb => 
                           mult_125_G3_FS_1_PG_int_0_4_0_port);
   U6520 : inv port map( inb => mult_125_G3_A1_17_port, outb => n5954);
   U6521 : inv port map( inb => mult_125_G3_A2_17_port, outb => n5955);
   U6522 : inv port map( inb => n5956, outb => 
                           mult_125_G3_FS_1_PG_int_0_4_1_port);
   U6523 : inv port map( inb => n5957, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_4_1_port);
   U6524 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_4_0_port, outb => 
                           n5958);
   U6525 : inv port map( inb => mult_125_G3_A1_18_port, outb => n5959);
   U6526 : inv port map( inb => mult_125_G3_A2_18_port, outb => n5960);
   U6527 : inv port map( inb => n5961, outb => 
                           mult_125_G3_FS_1_PG_int_0_4_2_port);
   U6528 : inv port map( inb => n5962, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_4_2_port);
   U6529 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_4_1_port, outb => 
                           n5963);
   U6530 : inv port map( inb => mult_125_G3_FS_1_C_1_4_1_port, outb => n5964);
   U6531 : inv port map( inb => mult_125_G3_FS_1_P_0_4_1_port, outb => n5965);
   U6532 : inv port map( inb => mult_125_G3_A1_19_port, outb => n5966);
   U6533 : inv port map( inb => mult_125_G3_A2_19_port, outb => n5967);
   U6534 : inv port map( inb => n5968, outb => 
                           mult_125_G3_FS_1_PG_int_0_4_3_port);
   U6535 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_4_2_port, outb => 
                           n5969);
   U6536 : inv port map( inb => mult_125_G3_FS_1_P_0_4_3_port, outb => n5970);
   U6537 : inv port map( inb => mult_125_G3_FS_1_C_1_4_2_port, outb => n5971);
   U6538 : inv port map( inb => mult_125_G3_FS_1_P_0_4_2_port, outb => n5972);
   U6539 : inv port map( inb => mult_125_G3_A1_20_port, outb => n5973);
   U6540 : inv port map( inb => mult_125_G3_A2_20_port, outb => n5974);
   U6541 : inv port map( inb => n5975, outb => 
                           mult_125_G3_FS_1_PG_int_0_5_0_port);
   U6542 : inv port map( inb => mult_125_G3_A1_21_port, outb => n5976);
   U6543 : inv port map( inb => mult_125_G3_A2_21_port, outb => n5977);
   U6544 : inv port map( inb => n5978, outb => 
                           mult_125_G3_FS_1_PG_int_0_5_1_port);
   U6545 : inv port map( inb => n5979, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_5_1_port);
   U6546 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_5_0_port, outb => 
                           n5980);
   U6547 : inv port map( inb => mult_125_G3_A1_22_port, outb => n5981);
   U6548 : inv port map( inb => mult_125_G3_A2_22_port, outb => n5982);
   U6549 : inv port map( inb => n5983, outb => 
                           mult_125_G3_FS_1_PG_int_0_5_2_port);
   U6550 : inv port map( inb => n5984, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_5_2_port);
   U6551 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_5_1_port, outb => 
                           n5985);
   U6552 : inv port map( inb => mult_125_G3_FS_1_C_1_5_1_port, outb => n5986);
   U6553 : inv port map( inb => mult_125_G3_FS_1_P_0_5_1_port, outb => n5987);
   U6554 : inv port map( inb => mult_125_G3_A1_23_port, outb => n5988);
   U6555 : inv port map( inb => mult_125_G3_A2_23_port, outb => n5989);
   U6556 : inv port map( inb => n5990, outb => 
                           mult_125_G3_FS_1_PG_int_0_5_3_port);
   U6557 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_5_2_port, outb => 
                           n5991);
   U6558 : inv port map( inb => mult_125_G3_FS_1_P_0_5_3_port, outb => n5992);
   U6559 : inv port map( inb => mult_125_G3_FS_1_C_1_5_2_port, outb => n5993);
   U6560 : inv port map( inb => mult_125_G3_FS_1_P_0_5_2_port, outb => n5994);
   U6561 : inv port map( inb => mult_125_G3_A1_24_port, outb => n5995);
   U6562 : inv port map( inb => mult_125_G3_A2_24_port, outb => n5996);
   U6563 : inv port map( inb => n5997, outb => 
                           mult_125_G3_FS_1_PG_int_0_6_0_port);
   U6564 : inv port map( inb => mult_125_G3_A1_25_port, outb => n5998);
   U6565 : inv port map( inb => mult_125_G3_A2_25_port, outb => n5999);
   U6566 : inv port map( inb => n6000, outb => 
                           mult_125_G3_FS_1_PG_int_0_6_1_port);
   U6567 : inv port map( inb => n6001, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_6_1_port);
   U6568 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_6_0_port, outb => 
                           n6002);
   U6569 : inv port map( inb => mult_125_G3_A1_26_port, outb => n6003);
   U6570 : inv port map( inb => mult_125_G3_A2_26_port, outb => n6004);
   U6571 : inv port map( inb => n6005, outb => 
                           mult_125_G3_FS_1_PG_int_0_6_2_port);
   U6572 : inv port map( inb => n6006, outb => 
                           mult_125_G3_FS_1_TEMP_P_0_6_2_port);
   U6573 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_6_1_port, outb => 
                           n6007);
   U6574 : inv port map( inb => mult_125_G3_FS_1_C_1_6_1_port, outb => n6008);
   U6575 : inv port map( inb => mult_125_G3_FS_1_P_0_6_1_port, outb => n6009);
   U6576 : inv port map( inb => mult_125_G3_A1_27_port, outb => n6010);
   U6577 : inv port map( inb => mult_125_G3_A2_27_port, outb => n6011);
   U6578 : inv port map( inb => n6012, outb => 
                           mult_125_G3_FS_1_PG_int_0_6_3_port);
   U6579 : inv port map( inb => mult_125_G3_FS_1_TEMP_G_0_6_2_port, outb => 
                           n6013);
   U6580 : inv port map( inb => mult_125_G3_FS_1_P_0_6_3_port, outb => n6014);
   U6581 : inv port map( inb => mult_125_G3_FS_1_C_1_6_2_port, outb => n6015);
   U6582 : inv port map( inb => mult_125_G3_FS_1_P_0_6_2_port, outb => n6016);
   U6583 : inv port map( inb => mult_125_G3_A1_28_port, outb => n6017);
   U6584 : inv port map( inb => mult_125_G3_A2_28_port, outb => n6018);
   U6585 : inv port map( inb => n6019, outb => 
                           mult_125_G3_FS_1_PG_int_0_7_0_port);
   U6586 : inv port map( inb => mult_125_G3_A1_29_port, outb => n6020);
   U6587 : inv port map( inb => mult_125_G3_A2_29_port, outb => n6021);
   U6588 : inv port map( inb => n6022, outb => 
                           mult_125_G3_FS_1_PG_int_0_7_1_port);
   U6589 : inv port map( inb => mult_125_G3_FS_1_C_1_7_0_port, outb => n6023);
   U6590 : inv port map( inb => mult_125_G3_FS_1_TEMP_P_0_7_0_port, outb => 
                           n6024);
   U6591 : inv port map( inb => mult_125_G3_FS_1_G_1_0_3_port, outb => n6025);
   U6592 : inv port map( inb => mult_125_G3_FS_1_C_1_4_0_port, outb => n6026);
   U6593 : inv port map( inb => mult_125_G3_FS_1_G_1_1_0_port, outb => n6028);
   U6594 : inv port map( inb => mult_125_G3_FS_1_C_1_5_0_port, outb => n6029);
   U6595 : inv port map( inb => mult_125_G3_FS_1_G_1_1_1_port, outb => n6031);
   U6596 : inv port map( inb => mult_125_G3_FS_1_C_1_6_0_port, outb => n6032);
   U6597 : inv port map( inb => mult_125_G3_FS_1_G_1_1_2_port, outb => n6034);
   U6598 : inv port map( inb => mult_125_G3_FS_1_G_2_0_0_port, outb => n6035);

end SYN_fir_rtl_arch;
