////////////////////////////////////////////////////////////////////////////////
// Module Name  : template_task_functions
// File name    : template_task_functions.sv
// Description  : Template for SystemVerilog Tasks and Functions
// Type         : 
// Limitations  : None
// Model Styles : 
// Author       : Varun Nagpal
// Revision|Date: 0.1 | 14/10/2020
////////////////////////////////////////////////////////////////////////////////